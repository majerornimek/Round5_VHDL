library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
use ieee.numeric_std.all;
-- use ieee.std_logic_arith.all;

library work;
use work.Round5_constants.all;

entity Unlift_Poly is 
	port (
		PolyA	: in q_bitsPoly(PolyDegree downto 0);
		clk 	: in std_logic;
		Start	: in std_logic;
		Done	: out std_logic;
		LongRes	: out q_bitsPoly(PolyDegree downto 0)
		-- ShortRes: out ShortPoly(PolyDegree downto 0)
	);
end entity;

architecture a1 of Unlift_Poly is
signal Long_tmp     : std_logic_vector(q_bits-1 downto 0);
signal counter	    : std_logic_vector(PolyDegreeLog2-1 downto 0);
signal PolyA_tmp    : q_bitsPoly(PolyDegree downto 0);
signal CycPoly_tmp  : q_bitsPoly(PolyDegree downto 0);
signal tmp_res	    : std_logic_vector(q_bits-1 downto 0);

signal ShortPolyTmp : p_bitsPoly(PolyDegree downto 0);

signal done_tmp     : std_logic;
begin

	

	
arithm: process(clk)
begin
	if clk'event and clk = '1' then
		if Start = '1' then
			if counter = 0 then
				tmp_res <= (others => '0');
			elsif counter = "00000000001" then
				tmp_res <= not PolyA(PolyDegree) + '1';
			else --if counter > 2 then
				tmp_res <= ( tmp_res - PolyA_tmp(PolyDegree));
			end if;
		else
			tmp_res <= (others => '0');
		end if;
	end if;
end process;


shift_poly: process(clk)
begin
	if clk'event and clk = '1' then
		if Start = '1' then
			if counter = 0 then
				PolyA_tmp <= PolyA;
			elsif counter < PolyDegree+1 then
				PolyA_tmp <= PolyA_tmp(PolyDegree-1 downto 0) & PolyA_tmp(PolyDegree);
			end if;
		end if;
	end if;
end process;

shift_cyc: process(clk)
begin
	if clk'event and clk = '1' then
		if Start = '1' then
			if counter = 0 then
			elsif counter = 1 then
			elsif counter < PolyDegree+3 then
				CycPoly_tmp <= CycPoly_tmp(PolyDegree-1 downto 0) & tmp_res;
			end if;
		else
			CycPoly_tmp <= (others =>(others=>'0'));
		end if;
	end if;
end process;
	
count: process(clk)
begin
	if clk'event and clk = '1' then
		if Start = '1' then
			if counter < PolyDegree+3 then
				counter <= counter + '1';
				done_tmp <= '0';
			else
				LongRes <= CycPoly_tmp;
				done_tmp <= '1';
			end if;
		else
			counter <= (others => '0');
			done_tmp <= '0';
		end if;
	end if;
end process;

Done <= done_tmp and start;
	
	
end a1;


-- architecture a2 of Unlift_Poly is
-- signal Long_tmp     : std_logic_vector(q_bits-1 downto 0);
-- signal input_pointer	    : std_logic_vector(PolyDegreeLog2-2 downto 0);
-- signal PolyA_tmp    : q_bitsPoly(PolyDegree downto 0);
-- signal CycPoly_tmp  : q_bitsPoly(PolyDegree downto 0);
-- signal tmp_res	    : std_logic_vector(q_bits-1 downto 0);

-- signal sub_element  : std_logic_vector(q_bits-1 downto 0);
-- signal sub_result   : std_logic_vector(q_bits-1 downto 0);
-- signal ShortPolyTmp : p_bitsPoly(PolyDegree downto 0);

-- signal done_tmp     : std_logic;
-- begin

-- process(clk)
-- begin
	-- if clk'event and clk = '1' then
		-- if Start = '1' then
			-- if input_pointer = 0 then
				-- sub_result <= (others => '0');
			-- elsif input_pointer = "00000000001" then
				-- sub_result <= not PolyA(PolyDegree) + '1';
			-- else --if counter > 2 then
				-- sub_result <= ( sub_result - sub_element);
			-- end if;
		-- else
			-- sub_result <= (others => '0');
		-- end if;
	-- end if;
-- end process;

	
	
-- count: process(clk)
-- begin
	-- if clk'event and clk = '1' then
		-- if Start = '1' then
			-- if input_pointer < PolyDegree+3 then
				-- input_pointer <= input_pointer + '1';
				-- done_tmp <= '0';
			-- else
				-- done_tmp <= '1';
			-- end if;
		-- else
			-- input_pointer <= (others => '0');
			-- done_tmp <= '0';
		-- end if;
	-- end if;
-- end process;

-- Done <= done_tmp and start;
	
----==========   InPUT Pointer  ================
-- process(clk)
-- begin
 -- if clk'event and clk = '1' then
     -- case input_pointer is

        -- when "0000000001" => 
-- sub_element <= PolyA(1018);
        -- when "0000000010" => 
-- sub_element <= PolyA(1017);
        -- when "0000000011" => 
-- sub_element <= PolyA(1016);
        -- when "0000000100" => 
-- sub_element <= PolyA(1015);
        -- when "0000000101" => 
-- sub_element <= PolyA(1014);
        -- when "0000000110" => 
-- sub_element <= PolyA(1013);
        -- when "0000000111" => 
-- sub_element <= PolyA(1012);
        -- when "0000001000" => 
-- sub_element <= PolyA(1011);
        -- when "0000001001" => 
-- sub_element <= PolyA(1010);
        -- when "0000001010" => 
-- sub_element <= PolyA(1009);
        -- when "0000001011" => 
-- sub_element <= PolyA(1008);
        -- when "0000001100" => 
-- sub_element <= PolyA(1007);
        -- when "0000001101" => 
-- sub_element <= PolyA(1006);
        -- when "0000001110" => 
-- sub_element <= PolyA(1005);
        -- when "0000001111" => 
-- sub_element <= PolyA(1004);
        -- when "0000010000" => 
-- sub_element <= PolyA(1003);
        -- when "0000010001" => 
-- sub_element <= PolyA(1002);
        -- when "0000010010" => 
-- sub_element <= PolyA(1001);
        -- when "0000010011" => 
-- sub_element <= PolyA(1000);
        -- when "0000010100" => 
-- sub_element <= PolyA(999);
        -- when "0000010101" => 
-- sub_element <= PolyA(998);
        -- when "0000010110" => 
-- sub_element <= PolyA(997);
        -- when "0000010111" => 
-- sub_element <= PolyA(996);
        -- when "0000011000" => 
-- sub_element <= PolyA(995);
        -- when "0000011001" => 
-- sub_element <= PolyA(994);
        -- when "0000011010" => 
-- sub_element <= PolyA(993);
        -- when "0000011011" => 
-- sub_element <= PolyA(992);
        -- when "0000011100" => 
-- sub_element <= PolyA(991);
        -- when "0000011101" => 
-- sub_element <= PolyA(990);
        -- when "0000011110" => 
-- sub_element <= PolyA(989);
        -- when "0000011111" => 
-- sub_element <= PolyA(988);
        -- when "0000100000" => 
-- sub_element <= PolyA(987);
        -- when "0000100001" => 
-- sub_element <= PolyA(986);
        -- when "0000100010" => 
-- sub_element <= PolyA(985);
        -- when "0000100011" => 
-- sub_element <= PolyA(984);
        -- when "0000100100" => 
-- sub_element <= PolyA(983);
        -- when "0000100101" => 
-- sub_element <= PolyA(982);
        -- when "0000100110" => 
-- sub_element <= PolyA(981);
        -- when "0000100111" => 
-- sub_element <= PolyA(980);
        -- when "0000101000" => 
-- sub_element <= PolyA(979);
        -- when "0000101001" => 
-- sub_element <= PolyA(978);
        -- when "0000101010" => 
-- sub_element <= PolyA(977);
        -- when "0000101011" => 
-- sub_element <= PolyA(976);
        -- when "0000101100" => 
-- sub_element <= PolyA(975);
        -- when "0000101101" => 
-- sub_element <= PolyA(974);
        -- when "0000101110" => 
-- sub_element <= PolyA(973);
        -- when "0000101111" => 
-- sub_element <= PolyA(972);
        -- when "0000110000" => 
-- sub_element <= PolyA(971);
        -- when "0000110001" => 
-- sub_element <= PolyA(970);
        -- when "0000110010" => 
-- sub_element <= PolyA(969);
        -- when "0000110011" => 
-- sub_element <= PolyA(968);
        -- when "0000110100" => 
-- sub_element <= PolyA(967);
        -- when "0000110101" => 
-- sub_element <= PolyA(966);
        -- when "0000110110" => 
-- sub_element <= PolyA(965);
        -- when "0000110111" => 
-- sub_element <= PolyA(964);
        -- when "0000111000" => 
-- sub_element <= PolyA(963);
        -- when "0000111001" => 
-- sub_element <= PolyA(962);
        -- when "0000111010" => 
-- sub_element <= PolyA(961);
        -- when "0000111011" => 
-- sub_element <= PolyA(960);
        -- when "0000111100" => 
-- sub_element <= PolyA(959);
        -- when "0000111101" => 
-- sub_element <= PolyA(958);
        -- when "0000111110" => 
-- sub_element <= PolyA(957);
        -- when "0000111111" => 
-- sub_element <= PolyA(956);
        -- when "0001000000" => 
-- sub_element <= PolyA(955);
        -- when "0001000001" => 
-- sub_element <= PolyA(954);
        -- when "0001000010" => 
-- sub_element <= PolyA(953);
        -- when "0001000011" => 
-- sub_element <= PolyA(952);
        -- when "0001000100" => 
-- sub_element <= PolyA(951);
        -- when "0001000101" => 
-- sub_element <= PolyA(950);
        -- when "0001000110" => 
-- sub_element <= PolyA(949);
        -- when "0001000111" => 
-- sub_element <= PolyA(948);
        -- when "0001001000" => 
-- sub_element <= PolyA(947);
        -- when "0001001001" => 
-- sub_element <= PolyA(946);
        -- when "0001001010" => 
-- sub_element <= PolyA(945);
        -- when "0001001011" => 
-- sub_element <= PolyA(944);
        -- when "0001001100" => 
-- sub_element <= PolyA(943);
        -- when "0001001101" => 
-- sub_element <= PolyA(942);
        -- when "0001001110" => 
-- sub_element <= PolyA(941);
        -- when "0001001111" => 
-- sub_element <= PolyA(940);
        -- when "0001010000" => 
-- sub_element <= PolyA(939);
        -- when "0001010001" => 
-- sub_element <= PolyA(938);
        -- when "0001010010" => 
-- sub_element <= PolyA(937);
        -- when "0001010011" => 
-- sub_element <= PolyA(936);
        -- when "0001010100" => 
-- sub_element <= PolyA(935);
        -- when "0001010101" => 
-- sub_element <= PolyA(934);
        -- when "0001010110" => 
-- sub_element <= PolyA(933);
        -- when "0001010111" => 
-- sub_element <= PolyA(932);
        -- when "0001011000" => 
-- sub_element <= PolyA(931);
        -- when "0001011001" => 
-- sub_element <= PolyA(930);
        -- when "0001011010" => 
-- sub_element <= PolyA(929);
        -- when "0001011011" => 
-- sub_element <= PolyA(928);
        -- when "0001011100" => 
-- sub_element <= PolyA(927);
        -- when "0001011101" => 
-- sub_element <= PolyA(926);
        -- when "0001011110" => 
-- sub_element <= PolyA(925);
        -- when "0001011111" => 
-- sub_element <= PolyA(924);
        -- when "0001100000" => 
-- sub_element <= PolyA(923);
        -- when "0001100001" => 
-- sub_element <= PolyA(922);
        -- when "0001100010" => 
-- sub_element <= PolyA(921);
        -- when "0001100011" => 
-- sub_element <= PolyA(920);
        -- when "0001100100" => 
-- sub_element <= PolyA(919);
        -- when "0001100101" => 
-- sub_element <= PolyA(918);
        -- when "0001100110" => 
-- sub_element <= PolyA(917);
        -- when "0001100111" => 
-- sub_element <= PolyA(916);
        -- when "0001101000" => 
-- sub_element <= PolyA(915);
        -- when "0001101001" => 
-- sub_element <= PolyA(914);
        -- when "0001101010" => 
-- sub_element <= PolyA(913);
        -- when "0001101011" => 
-- sub_element <= PolyA(912);
        -- when "0001101100" => 
-- sub_element <= PolyA(911);
        -- when "0001101101" => 
-- sub_element <= PolyA(910);
        -- when "0001101110" => 
-- sub_element <= PolyA(909);
        -- when "0001101111" => 
-- sub_element <= PolyA(908);
        -- when "0001110000" => 
-- sub_element <= PolyA(907);
        -- when "0001110001" => 
-- sub_element <= PolyA(906);
        -- when "0001110010" => 
-- sub_element <= PolyA(905);
        -- when "0001110011" => 
-- sub_element <= PolyA(904);
        -- when "0001110100" => 
-- sub_element <= PolyA(903);
        -- when "0001110101" => 
-- sub_element <= PolyA(902);
        -- when "0001110110" => 
-- sub_element <= PolyA(901);
        -- when "0001110111" => 
-- sub_element <= PolyA(900);
        -- when "0001111000" => 
-- sub_element <= PolyA(899);
        -- when "0001111001" => 
-- sub_element <= PolyA(898);
        -- when "0001111010" => 
-- sub_element <= PolyA(897);
        -- when "0001111011" => 
-- sub_element <= PolyA(896);
        -- when "0001111100" => 
-- sub_element <= PolyA(895);
        -- when "0001111101" => 
-- sub_element <= PolyA(894);
        -- when "0001111110" => 
-- sub_element <= PolyA(893);
        -- when "0001111111" => 
-- sub_element <= PolyA(892);
        -- when "0010000000" => 
-- sub_element <= PolyA(891);
        -- when "0010000001" => 
-- sub_element <= PolyA(890);
        -- when "0010000010" => 
-- sub_element <= PolyA(889);
        -- when "0010000011" => 
-- sub_element <= PolyA(888);
        -- when "0010000100" => 
-- sub_element <= PolyA(887);
        -- when "0010000101" => 
-- sub_element <= PolyA(886);
        -- when "0010000110" => 
-- sub_element <= PolyA(885);
        -- when "0010000111" => 
-- sub_element <= PolyA(884);
        -- when "0010001000" => 
-- sub_element <= PolyA(883);
        -- when "0010001001" => 
-- sub_element <= PolyA(882);
        -- when "0010001010" => 
-- sub_element <= PolyA(881);
        -- when "0010001011" => 
-- sub_element <= PolyA(880);
        -- when "0010001100" => 
-- sub_element <= PolyA(879);
        -- when "0010001101" => 
-- sub_element <= PolyA(878);
        -- when "0010001110" => 
-- sub_element <= PolyA(877);
        -- when "0010001111" => 
-- sub_element <= PolyA(876);
        -- when "0010010000" => 
-- sub_element <= PolyA(875);
        -- when "0010010001" => 
-- sub_element <= PolyA(874);
        -- when "0010010010" => 
-- sub_element <= PolyA(873);
        -- when "0010010011" => 
-- sub_element <= PolyA(872);
        -- when "0010010100" => 
-- sub_element <= PolyA(871);
        -- when "0010010101" => 
-- sub_element <= PolyA(870);
        -- when "0010010110" => 
-- sub_element <= PolyA(869);
        -- when "0010010111" => 
-- sub_element <= PolyA(868);
        -- when "0010011000" => 
-- sub_element <= PolyA(867);
        -- when "0010011001" => 
-- sub_element <= PolyA(866);
        -- when "0010011010" => 
-- sub_element <= PolyA(865);
        -- when "0010011011" => 
-- sub_element <= PolyA(864);
        -- when "0010011100" => 
-- sub_element <= PolyA(863);
        -- when "0010011101" => 
-- sub_element <= PolyA(862);
        -- when "0010011110" => 
-- sub_element <= PolyA(861);
        -- when "0010011111" => 
-- sub_element <= PolyA(860);
        -- when "0010100000" => 
-- sub_element <= PolyA(859);
        -- when "0010100001" => 
-- sub_element <= PolyA(858);
        -- when "0010100010" => 
-- sub_element <= PolyA(857);
        -- when "0010100011" => 
-- sub_element <= PolyA(856);
        -- when "0010100100" => 
-- sub_element <= PolyA(855);
        -- when "0010100101" => 
-- sub_element <= PolyA(854);
        -- when "0010100110" => 
-- sub_element <= PolyA(853);
        -- when "0010100111" => 
-- sub_element <= PolyA(852);
        -- when "0010101000" => 
-- sub_element <= PolyA(851);
        -- when "0010101001" => 
-- sub_element <= PolyA(850);
        -- when "0010101010" => 
-- sub_element <= PolyA(849);
        -- when "0010101011" => 
-- sub_element <= PolyA(848);
        -- when "0010101100" => 
-- sub_element <= PolyA(847);
        -- when "0010101101" => 
-- sub_element <= PolyA(846);
        -- when "0010101110" => 
-- sub_element <= PolyA(845);
        -- when "0010101111" => 
-- sub_element <= PolyA(844);
        -- when "0010110000" => 
-- sub_element <= PolyA(843);
        -- when "0010110001" => 
-- sub_element <= PolyA(842);
        -- when "0010110010" => 
-- sub_element <= PolyA(841);
        -- when "0010110011" => 
-- sub_element <= PolyA(840);
        -- when "0010110100" => 
-- sub_element <= PolyA(839);
        -- when "0010110101" => 
-- sub_element <= PolyA(838);
        -- when "0010110110" => 
-- sub_element <= PolyA(837);
        -- when "0010110111" => 
-- sub_element <= PolyA(836);
        -- when "0010111000" => 
-- sub_element <= PolyA(835);
        -- when "0010111001" => 
-- sub_element <= PolyA(834);
        -- when "0010111010" => 
-- sub_element <= PolyA(833);
        -- when "0010111011" => 
-- sub_element <= PolyA(832);
        -- when "0010111100" => 
-- sub_element <= PolyA(831);
        -- when "0010111101" => 
-- sub_element <= PolyA(830);
        -- when "0010111110" => 
-- sub_element <= PolyA(829);
        -- when "0010111111" => 
-- sub_element <= PolyA(828);
        -- when "0011000000" => 
-- sub_element <= PolyA(827);
        -- when "0011000001" => 
-- sub_element <= PolyA(826);
        -- when "0011000010" => 
-- sub_element <= PolyA(825);
        -- when "0011000011" => 
-- sub_element <= PolyA(824);
        -- when "0011000100" => 
-- sub_element <= PolyA(823);
        -- when "0011000101" => 
-- sub_element <= PolyA(822);
        -- when "0011000110" => 
-- sub_element <= PolyA(821);
        -- when "0011000111" => 
-- sub_element <= PolyA(820);
        -- when "0011001000" => 
-- sub_element <= PolyA(819);
        -- when "0011001001" => 
-- sub_element <= PolyA(818);
        -- when "0011001010" => 
-- sub_element <= PolyA(817);
        -- when "0011001011" => 
-- sub_element <= PolyA(816);
        -- when "0011001100" => 
-- sub_element <= PolyA(815);
        -- when "0011001101" => 
-- sub_element <= PolyA(814);
        -- when "0011001110" => 
-- sub_element <= PolyA(813);
        -- when "0011001111" => 
-- sub_element <= PolyA(812);
        -- when "0011010000" => 
-- sub_element <= PolyA(811);
        -- when "0011010001" => 
-- sub_element <= PolyA(810);
        -- when "0011010010" => 
-- sub_element <= PolyA(809);
        -- when "0011010011" => 
-- sub_element <= PolyA(808);
        -- when "0011010100" => 
-- sub_element <= PolyA(807);
        -- when "0011010101" => 
-- sub_element <= PolyA(806);
        -- when "0011010110" => 
-- sub_element <= PolyA(805);
        -- when "0011010111" => 
-- sub_element <= PolyA(804);
        -- when "0011011000" => 
-- sub_element <= PolyA(803);
        -- when "0011011001" => 
-- sub_element <= PolyA(802);
        -- when "0011011010" => 
-- sub_element <= PolyA(801);
        -- when "0011011011" => 
-- sub_element <= PolyA(800);
        -- when "0011011100" => 
-- sub_element <= PolyA(799);
        -- when "0011011101" => 
-- sub_element <= PolyA(798);
        -- when "0011011110" => 
-- sub_element <= PolyA(797);
        -- when "0011011111" => 
-- sub_element <= PolyA(796);
        -- when "0011100000" => 
-- sub_element <= PolyA(795);
        -- when "0011100001" => 
-- sub_element <= PolyA(794);
        -- when "0011100010" => 
-- sub_element <= PolyA(793);
        -- when "0011100011" => 
-- sub_element <= PolyA(792);
        -- when "0011100100" => 
-- sub_element <= PolyA(791);
        -- when "0011100101" => 
-- sub_element <= PolyA(790);
        -- when "0011100110" => 
-- sub_element <= PolyA(789);
        -- when "0011100111" => 
-- sub_element <= PolyA(788);
        -- when "0011101000" => 
-- sub_element <= PolyA(787);
        -- when "0011101001" => 
-- sub_element <= PolyA(786);
        -- when "0011101010" => 
-- sub_element <= PolyA(785);
        -- when "0011101011" => 
-- sub_element <= PolyA(784);
        -- when "0011101100" => 
-- sub_element <= PolyA(783);
        -- when "0011101101" => 
-- sub_element <= PolyA(782);
        -- when "0011101110" => 
-- sub_element <= PolyA(781);
        -- when "0011101111" => 
-- sub_element <= PolyA(780);
        -- when "0011110000" => 
-- sub_element <= PolyA(779);
        -- when "0011110001" => 
-- sub_element <= PolyA(778);
        -- when "0011110010" => 
-- sub_element <= PolyA(777);
        -- when "0011110011" => 
-- sub_element <= PolyA(776);
        -- when "0011110100" => 
-- sub_element <= PolyA(775);
        -- when "0011110101" => 
-- sub_element <= PolyA(774);
        -- when "0011110110" => 
-- sub_element <= PolyA(773);
        -- when "0011110111" => 
-- sub_element <= PolyA(772);
        -- when "0011111000" => 
-- sub_element <= PolyA(771);
        -- when "0011111001" => 
-- sub_element <= PolyA(770);
        -- when "0011111010" => 
-- sub_element <= PolyA(769);
        -- when "0011111011" => 
-- sub_element <= PolyA(768);
        -- when "0011111100" => 
-- sub_element <= PolyA(767);
        -- when "0011111101" => 
-- sub_element <= PolyA(766);
        -- when "0011111110" => 
-- sub_element <= PolyA(765);
        -- when "0011111111" => 
-- sub_element <= PolyA(764);
        -- when "0100000000" => 
-- sub_element <= PolyA(763);
        -- when "0100000001" => 
-- sub_element <= PolyA(762);
        -- when "0100000010" => 
-- sub_element <= PolyA(761);
        -- when "0100000011" => 
-- sub_element <= PolyA(760);
        -- when "0100000100" => 
-- sub_element <= PolyA(759);
        -- when "0100000101" => 
-- sub_element <= PolyA(758);
        -- when "0100000110" => 
-- sub_element <= PolyA(757);
        -- when "0100000111" => 
-- sub_element <= PolyA(756);
        -- when "0100001000" => 
-- sub_element <= PolyA(755);
        -- when "0100001001" => 
-- sub_element <= PolyA(754);
        -- when "0100001010" => 
-- sub_element <= PolyA(753);
        -- when "0100001011" => 
-- sub_element <= PolyA(752);
        -- when "0100001100" => 
-- sub_element <= PolyA(751);
        -- when "0100001101" => 
-- sub_element <= PolyA(750);
        -- when "0100001110" => 
-- sub_element <= PolyA(749);
        -- when "0100001111" => 
-- sub_element <= PolyA(748);
        -- when "0100010000" => 
-- sub_element <= PolyA(747);
        -- when "0100010001" => 
-- sub_element <= PolyA(746);
        -- when "0100010010" => 
-- sub_element <= PolyA(745);
        -- when "0100010011" => 
-- sub_element <= PolyA(744);
        -- when "0100010100" => 
-- sub_element <= PolyA(743);
        -- when "0100010101" => 
-- sub_element <= PolyA(742);
        -- when "0100010110" => 
-- sub_element <= PolyA(741);
        -- when "0100010111" => 
-- sub_element <= PolyA(740);
        -- when "0100011000" => 
-- sub_element <= PolyA(739);
        -- when "0100011001" => 
-- sub_element <= PolyA(738);
        -- when "0100011010" => 
-- sub_element <= PolyA(737);
        -- when "0100011011" => 
-- sub_element <= PolyA(736);
        -- when "0100011100" => 
-- sub_element <= PolyA(735);
        -- when "0100011101" => 
-- sub_element <= PolyA(734);
        -- when "0100011110" => 
-- sub_element <= PolyA(733);
        -- when "0100011111" => 
-- sub_element <= PolyA(732);
        -- when "0100100000" => 
-- sub_element <= PolyA(731);
        -- when "0100100001" => 
-- sub_element <= PolyA(730);
        -- when "0100100010" => 
-- sub_element <= PolyA(729);
        -- when "0100100011" => 
-- sub_element <= PolyA(728);
        -- when "0100100100" => 
-- sub_element <= PolyA(727);
        -- when "0100100101" => 
-- sub_element <= PolyA(726);
        -- when "0100100110" => 
-- sub_element <= PolyA(725);
        -- when "0100100111" => 
-- sub_element <= PolyA(724);
        -- when "0100101000" => 
-- sub_element <= PolyA(723);
        -- when "0100101001" => 
-- sub_element <= PolyA(722);
        -- when "0100101010" => 
-- sub_element <= PolyA(721);
        -- when "0100101011" => 
-- sub_element <= PolyA(720);
        -- when "0100101100" => 
-- sub_element <= PolyA(719);
        -- when "0100101101" => 
-- sub_element <= PolyA(718);
        -- when "0100101110" => 
-- sub_element <= PolyA(717);
        -- when "0100101111" => 
-- sub_element <= PolyA(716);
        -- when "0100110000" => 
-- sub_element <= PolyA(715);
        -- when "0100110001" => 
-- sub_element <= PolyA(714);
        -- when "0100110010" => 
-- sub_element <= PolyA(713);
        -- when "0100110011" => 
-- sub_element <= PolyA(712);
        -- when "0100110100" => 
-- sub_element <= PolyA(711);
        -- when "0100110101" => 
-- sub_element <= PolyA(710);
        -- when "0100110110" => 
-- sub_element <= PolyA(709);
        -- when "0100110111" => 
-- sub_element <= PolyA(708);
        -- when "0100111000" => 
-- sub_element <= PolyA(707);
        -- when "0100111001" => 
-- sub_element <= PolyA(706);
        -- when "0100111010" => 
-- sub_element <= PolyA(705);
        -- when "0100111011" => 
-- sub_element <= PolyA(704);
        -- when "0100111100" => 
-- sub_element <= PolyA(703);
        -- when "0100111101" => 
-- sub_element <= PolyA(702);
        -- when "0100111110" => 
-- sub_element <= PolyA(701);
        -- when "0100111111" => 
-- sub_element <= PolyA(700);
        -- when "0101000000" => 
-- sub_element <= PolyA(699);
        -- when "0101000001" => 
-- sub_element <= PolyA(698);
        -- when "0101000010" => 
-- sub_element <= PolyA(697);
        -- when "0101000011" => 
-- sub_element <= PolyA(696);
        -- when "0101000100" => 
-- sub_element <= PolyA(695);
        -- when "0101000101" => 
-- sub_element <= PolyA(694);
        -- when "0101000110" => 
-- sub_element <= PolyA(693);
        -- when "0101000111" => 
-- sub_element <= PolyA(692);
        -- when "0101001000" => 
-- sub_element <= PolyA(691);
        -- when "0101001001" => 
-- sub_element <= PolyA(690);
        -- when "0101001010" => 
-- sub_element <= PolyA(689);
        -- when "0101001011" => 
-- sub_element <= PolyA(688);
        -- when "0101001100" => 
-- sub_element <= PolyA(687);
        -- when "0101001101" => 
-- sub_element <= PolyA(686);
        -- when "0101001110" => 
-- sub_element <= PolyA(685);
        -- when "0101001111" => 
-- sub_element <= PolyA(684);
        -- when "0101010000" => 
-- sub_element <= PolyA(683);
        -- when "0101010001" => 
-- sub_element <= PolyA(682);
        -- when "0101010010" => 
-- sub_element <= PolyA(681);
        -- when "0101010011" => 
-- sub_element <= PolyA(680);
        -- when "0101010100" => 
-- sub_element <= PolyA(679);
        -- when "0101010101" => 
-- sub_element <= PolyA(678);
        -- when "0101010110" => 
-- sub_element <= PolyA(677);
        -- when "0101010111" => 
-- sub_element <= PolyA(676);
        -- when "0101011000" => 
-- sub_element <= PolyA(675);
        -- when "0101011001" => 
-- sub_element <= PolyA(674);
        -- when "0101011010" => 
-- sub_element <= PolyA(673);
        -- when "0101011011" => 
-- sub_element <= PolyA(672);
        -- when "0101011100" => 
-- sub_element <= PolyA(671);
        -- when "0101011101" => 
-- sub_element <= PolyA(670);
        -- when "0101011110" => 
-- sub_element <= PolyA(669);
        -- when "0101011111" => 
-- sub_element <= PolyA(668);
        -- when "0101100000" => 
-- sub_element <= PolyA(667);
        -- when "0101100001" => 
-- sub_element <= PolyA(666);
        -- when "0101100010" => 
-- sub_element <= PolyA(665);
        -- when "0101100011" => 
-- sub_element <= PolyA(664);
        -- when "0101100100" => 
-- sub_element <= PolyA(663);
        -- when "0101100101" => 
-- sub_element <= PolyA(662);
        -- when "0101100110" => 
-- sub_element <= PolyA(661);
        -- when "0101100111" => 
-- sub_element <= PolyA(660);
        -- when "0101101000" => 
-- sub_element <= PolyA(659);
        -- when "0101101001" => 
-- sub_element <= PolyA(658);
        -- when "0101101010" => 
-- sub_element <= PolyA(657);
        -- when "0101101011" => 
-- sub_element <= PolyA(656);
        -- when "0101101100" => 
-- sub_element <= PolyA(655);
        -- when "0101101101" => 
-- sub_element <= PolyA(654);
        -- when "0101101110" => 
-- sub_element <= PolyA(653);
        -- when "0101101111" => 
-- sub_element <= PolyA(652);
        -- when "0101110000" => 
-- sub_element <= PolyA(651);
        -- when "0101110001" => 
-- sub_element <= PolyA(650);
        -- when "0101110010" => 
-- sub_element <= PolyA(649);
        -- when "0101110011" => 
-- sub_element <= PolyA(648);
        -- when "0101110100" => 
-- sub_element <= PolyA(647);
        -- when "0101110101" => 
-- sub_element <= PolyA(646);
        -- when "0101110110" => 
-- sub_element <= PolyA(645);
        -- when "0101110111" => 
-- sub_element <= PolyA(644);
        -- when "0101111000" => 
-- sub_element <= PolyA(643);
        -- when "0101111001" => 
-- sub_element <= PolyA(642);
        -- when "0101111010" => 
-- sub_element <= PolyA(641);
        -- when "0101111011" => 
-- sub_element <= PolyA(640);
        -- when "0101111100" => 
-- sub_element <= PolyA(639);
        -- when "0101111101" => 
-- sub_element <= PolyA(638);
        -- when "0101111110" => 
-- sub_element <= PolyA(637);
        -- when "0101111111" => 
-- sub_element <= PolyA(636);
        -- when "0110000000" => 
-- sub_element <= PolyA(635);
        -- when "0110000001" => 
-- sub_element <= PolyA(634);
        -- when "0110000010" => 
-- sub_element <= PolyA(633);
        -- when "0110000011" => 
-- sub_element <= PolyA(632);
        -- when "0110000100" => 
-- sub_element <= PolyA(631);
        -- when "0110000101" => 
-- sub_element <= PolyA(630);
        -- when "0110000110" => 
-- sub_element <= PolyA(629);
        -- when "0110000111" => 
-- sub_element <= PolyA(628);
        -- when "0110001000" => 
-- sub_element <= PolyA(627);
        -- when "0110001001" => 
-- sub_element <= PolyA(626);
        -- when "0110001010" => 
-- sub_element <= PolyA(625);
        -- when "0110001011" => 
-- sub_element <= PolyA(624);
        -- when "0110001100" => 
-- sub_element <= PolyA(623);
        -- when "0110001101" => 
-- sub_element <= PolyA(622);
        -- when "0110001110" => 
-- sub_element <= PolyA(621);
        -- when "0110001111" => 
-- sub_element <= PolyA(620);
        -- when "0110010000" => 
-- sub_element <= PolyA(619);
        -- when "0110010001" => 
-- sub_element <= PolyA(618);
        -- when "0110010010" => 
-- sub_element <= PolyA(617);
        -- when "0110010011" => 
-- sub_element <= PolyA(616);
        -- when "0110010100" => 
-- sub_element <= PolyA(615);
        -- when "0110010101" => 
-- sub_element <= PolyA(614);
        -- when "0110010110" => 
-- sub_element <= PolyA(613);
        -- when "0110010111" => 
-- sub_element <= PolyA(612);
        -- when "0110011000" => 
-- sub_element <= PolyA(611);
        -- when "0110011001" => 
-- sub_element <= PolyA(610);
        -- when "0110011010" => 
-- sub_element <= PolyA(609);
        -- when "0110011011" => 
-- sub_element <= PolyA(608);
        -- when "0110011100" => 
-- sub_element <= PolyA(607);
        -- when "0110011101" => 
-- sub_element <= PolyA(606);
        -- when "0110011110" => 
-- sub_element <= PolyA(605);
        -- when "0110011111" => 
-- sub_element <= PolyA(604);
        -- when "0110100000" => 
-- sub_element <= PolyA(603);
        -- when "0110100001" => 
-- sub_element <= PolyA(602);
        -- when "0110100010" => 
-- sub_element <= PolyA(601);
        -- when "0110100011" => 
-- sub_element <= PolyA(600);
        -- when "0110100100" => 
-- sub_element <= PolyA(599);
        -- when "0110100101" => 
-- sub_element <= PolyA(598);
        -- when "0110100110" => 
-- sub_element <= PolyA(597);
        -- when "0110100111" => 
-- sub_element <= PolyA(596);
        -- when "0110101000" => 
-- sub_element <= PolyA(595);
        -- when "0110101001" => 
-- sub_element <= PolyA(594);
        -- when "0110101010" => 
-- sub_element <= PolyA(593);
        -- when "0110101011" => 
-- sub_element <= PolyA(592);
        -- when "0110101100" => 
-- sub_element <= PolyA(591);
        -- when "0110101101" => 
-- sub_element <= PolyA(590);
        -- when "0110101110" => 
-- sub_element <= PolyA(589);
        -- when "0110101111" => 
-- sub_element <= PolyA(588);
        -- when "0110110000" => 
-- sub_element <= PolyA(587);
        -- when "0110110001" => 
-- sub_element <= PolyA(586);
        -- when "0110110010" => 
-- sub_element <= PolyA(585);
        -- when "0110110011" => 
-- sub_element <= PolyA(584);
        -- when "0110110100" => 
-- sub_element <= PolyA(583);
        -- when "0110110101" => 
-- sub_element <= PolyA(582);
        -- when "0110110110" => 
-- sub_element <= PolyA(581);
        -- when "0110110111" => 
-- sub_element <= PolyA(580);
        -- when "0110111000" => 
-- sub_element <= PolyA(579);
        -- when "0110111001" => 
-- sub_element <= PolyA(578);
        -- when "0110111010" => 
-- sub_element <= PolyA(577);
        -- when "0110111011" => 
-- sub_element <= PolyA(576);
        -- when "0110111100" => 
-- sub_element <= PolyA(575);
        -- when "0110111101" => 
-- sub_element <= PolyA(574);
        -- when "0110111110" => 
-- sub_element <= PolyA(573);
        -- when "0110111111" => 
-- sub_element <= PolyA(572);
        -- when "0111000000" => 
-- sub_element <= PolyA(571);
        -- when "0111000001" => 
-- sub_element <= PolyA(570);
        -- when "0111000010" => 
-- sub_element <= PolyA(569);
        -- when "0111000011" => 
-- sub_element <= PolyA(568);
        -- when "0111000100" => 
-- sub_element <= PolyA(567);
        -- when "0111000101" => 
-- sub_element <= PolyA(566);
        -- when "0111000110" => 
-- sub_element <= PolyA(565);
        -- when "0111000111" => 
-- sub_element <= PolyA(564);
        -- when "0111001000" => 
-- sub_element <= PolyA(563);
        -- when "0111001001" => 
-- sub_element <= PolyA(562);
        -- when "0111001010" => 
-- sub_element <= PolyA(561);
        -- when "0111001011" => 
-- sub_element <= PolyA(560);
        -- when "0111001100" => 
-- sub_element <= PolyA(559);
        -- when "0111001101" => 
-- sub_element <= PolyA(558);
        -- when "0111001110" => 
-- sub_element <= PolyA(557);
        -- when "0111001111" => 
-- sub_element <= PolyA(556);
        -- when "0111010000" => 
-- sub_element <= PolyA(555);
        -- when "0111010001" => 
-- sub_element <= PolyA(554);
        -- when "0111010010" => 
-- sub_element <= PolyA(553);
        -- when "0111010011" => 
-- sub_element <= PolyA(552);
        -- when "0111010100" => 
-- sub_element <= PolyA(551);
        -- when "0111010101" => 
-- sub_element <= PolyA(550);
        -- when "0111010110" => 
-- sub_element <= PolyA(549);
        -- when "0111010111" => 
-- sub_element <= PolyA(548);
        -- when "0111011000" => 
-- sub_element <= PolyA(547);
        -- when "0111011001" => 
-- sub_element <= PolyA(546);
        -- when "0111011010" => 
-- sub_element <= PolyA(545);
        -- when "0111011011" => 
-- sub_element <= PolyA(544);
        -- when "0111011100" => 
-- sub_element <= PolyA(543);
        -- when "0111011101" => 
-- sub_element <= PolyA(542);
        -- when "0111011110" => 
-- sub_element <= PolyA(541);
        -- when "0111011111" => 
-- sub_element <= PolyA(540);
        -- when "0111100000" => 
-- sub_element <= PolyA(539);
        -- when "0111100001" => 
-- sub_element <= PolyA(538);
        -- when "0111100010" => 
-- sub_element <= PolyA(537);
        -- when "0111100011" => 
-- sub_element <= PolyA(536);
        -- when "0111100100" => 
-- sub_element <= PolyA(535);
        -- when "0111100101" => 
-- sub_element <= PolyA(534);
        -- when "0111100110" => 
-- sub_element <= PolyA(533);
        -- when "0111100111" => 
-- sub_element <= PolyA(532);
        -- when "0111101000" => 
-- sub_element <= PolyA(531);
        -- when "0111101001" => 
-- sub_element <= PolyA(530);
        -- when "0111101010" => 
-- sub_element <= PolyA(529);
        -- when "0111101011" => 
-- sub_element <= PolyA(528);
        -- when "0111101100" => 
-- sub_element <= PolyA(527);
        -- when "0111101101" => 
-- sub_element <= PolyA(526);
        -- when "0111101110" => 
-- sub_element <= PolyA(525);
        -- when "0111101111" => 
-- sub_element <= PolyA(524);
        -- when "0111110000" => 
-- sub_element <= PolyA(523);
        -- when "0111110001" => 
-- sub_element <= PolyA(522);
        -- when "0111110010" => 
-- sub_element <= PolyA(521);
        -- when "0111110011" => 
-- sub_element <= PolyA(520);
        -- when "0111110100" => 
-- sub_element <= PolyA(519);
        -- when "0111110101" => 
-- sub_element <= PolyA(518);
        -- when "0111110110" => 
-- sub_element <= PolyA(517);
        -- when "0111110111" => 
-- sub_element <= PolyA(516);
        -- when "0111111000" => 
-- sub_element <= PolyA(515);
        -- when "0111111001" => 
-- sub_element <= PolyA(514);
        -- when "0111111010" => 
-- sub_element <= PolyA(513);
        -- when "0111111011" => 
-- sub_element <= PolyA(512);
        -- when "0111111100" => 
-- sub_element <= PolyA(511);
        -- when "0111111101" => 
-- sub_element <= PolyA(510);
        -- when "0111111110" => 
-- sub_element <= PolyA(509);
        -- when "0111111111" => 
-- sub_element <= PolyA(508);
        -- when "1000000000" => 
-- sub_element <= PolyA(507);
        -- when "1000000001" => 
-- sub_element <= PolyA(506);
        -- when "1000000010" => 
-- sub_element <= PolyA(505);
        -- when "1000000011" => 
-- sub_element <= PolyA(504);
        -- when "1000000100" => 
-- sub_element <= PolyA(503);
        -- when "1000000101" => 
-- sub_element <= PolyA(502);
        -- when "1000000110" => 
-- sub_element <= PolyA(501);
        -- when "1000000111" => 
-- sub_element <= PolyA(500);
        -- when "1000001000" => 
-- sub_element <= PolyA(499);
        -- when "1000001001" => 
-- sub_element <= PolyA(498);
        -- when "1000001010" => 
-- sub_element <= PolyA(497);
        -- when "1000001011" => 
-- sub_element <= PolyA(496);
        -- when "1000001100" => 
-- sub_element <= PolyA(495);
        -- when "1000001101" => 
-- sub_element <= PolyA(494);
        -- when "1000001110" => 
-- sub_element <= PolyA(493);
        -- when "1000001111" => 
-- sub_element <= PolyA(492);
        -- when "1000010000" => 
-- sub_element <= PolyA(491);
        -- when "1000010001" => 
-- sub_element <= PolyA(490);
        -- when "1000010010" => 
-- sub_element <= PolyA(489);
        -- when "1000010011" => 
-- sub_element <= PolyA(488);
        -- when "1000010100" => 
-- sub_element <= PolyA(487);
        -- when "1000010101" => 
-- sub_element <= PolyA(486);
        -- when "1000010110" => 
-- sub_element <= PolyA(485);
        -- when "1000010111" => 
-- sub_element <= PolyA(484);
        -- when "1000011000" => 
-- sub_element <= PolyA(483);
        -- when "1000011001" => 
-- sub_element <= PolyA(482);
        -- when "1000011010" => 
-- sub_element <= PolyA(481);
        -- when "1000011011" => 
-- sub_element <= PolyA(480);
        -- when "1000011100" => 
-- sub_element <= PolyA(479);
        -- when "1000011101" => 
-- sub_element <= PolyA(478);
        -- when "1000011110" => 
-- sub_element <= PolyA(477);
        -- when "1000011111" => 
-- sub_element <= PolyA(476);
        -- when "1000100000" => 
-- sub_element <= PolyA(475);
        -- when "1000100001" => 
-- sub_element <= PolyA(474);
        -- when "1000100010" => 
-- sub_element <= PolyA(473);
        -- when "1000100011" => 
-- sub_element <= PolyA(472);
        -- when "1000100100" => 
-- sub_element <= PolyA(471);
        -- when "1000100101" => 
-- sub_element <= PolyA(470);
        -- when "1000100110" => 
-- sub_element <= PolyA(469);
        -- when "1000100111" => 
-- sub_element <= PolyA(468);
        -- when "1000101000" => 
-- sub_element <= PolyA(467);
        -- when "1000101001" => 
-- sub_element <= PolyA(466);
        -- when "1000101010" => 
-- sub_element <= PolyA(465);
        -- when "1000101011" => 
-- sub_element <= PolyA(464);
        -- when "1000101100" => 
-- sub_element <= PolyA(463);
        -- when "1000101101" => 
-- sub_element <= PolyA(462);
        -- when "1000101110" => 
-- sub_element <= PolyA(461);
        -- when "1000101111" => 
-- sub_element <= PolyA(460);
        -- when "1000110000" => 
-- sub_element <= PolyA(459);
        -- when "1000110001" => 
-- sub_element <= PolyA(458);
        -- when "1000110010" => 
-- sub_element <= PolyA(457);
        -- when "1000110011" => 
-- sub_element <= PolyA(456);
        -- when "1000110100" => 
-- sub_element <= PolyA(455);
        -- when "1000110101" => 
-- sub_element <= PolyA(454);
        -- when "1000110110" => 
-- sub_element <= PolyA(453);
        -- when "1000110111" => 
-- sub_element <= PolyA(452);
        -- when "1000111000" => 
-- sub_element <= PolyA(451);
        -- when "1000111001" => 
-- sub_element <= PolyA(450);
        -- when "1000111010" => 
-- sub_element <= PolyA(449);
        -- when "1000111011" => 
-- sub_element <= PolyA(448);
        -- when "1000111100" => 
-- sub_element <= PolyA(447);
        -- when "1000111101" => 
-- sub_element <= PolyA(446);
        -- when "1000111110" => 
-- sub_element <= PolyA(445);
        -- when "1000111111" => 
-- sub_element <= PolyA(444);
        -- when "1001000000" => 
-- sub_element <= PolyA(443);
        -- when "1001000001" => 
-- sub_element <= PolyA(442);
        -- when "1001000010" => 
-- sub_element <= PolyA(441);
        -- when "1001000011" => 
-- sub_element <= PolyA(440);
        -- when "1001000100" => 
-- sub_element <= PolyA(439);
        -- when "1001000101" => 
-- sub_element <= PolyA(438);
        -- when "1001000110" => 
-- sub_element <= PolyA(437);
        -- when "1001000111" => 
-- sub_element <= PolyA(436);
        -- when "1001001000" => 
-- sub_element <= PolyA(435);
        -- when "1001001001" => 
-- sub_element <= PolyA(434);
        -- when "1001001010" => 
-- sub_element <= PolyA(433);
        -- when "1001001011" => 
-- sub_element <= PolyA(432);
        -- when "1001001100" => 
-- sub_element <= PolyA(431);
        -- when "1001001101" => 
-- sub_element <= PolyA(430);
        -- when "1001001110" => 
-- sub_element <= PolyA(429);
        -- when "1001001111" => 
-- sub_element <= PolyA(428);
        -- when "1001010000" => 
-- sub_element <= PolyA(427);
        -- when "1001010001" => 
-- sub_element <= PolyA(426);
        -- when "1001010010" => 
-- sub_element <= PolyA(425);
        -- when "1001010011" => 
-- sub_element <= PolyA(424);
        -- when "1001010100" => 
-- sub_element <= PolyA(423);
        -- when "1001010101" => 
-- sub_element <= PolyA(422);
        -- when "1001010110" => 
-- sub_element <= PolyA(421);
        -- when "1001010111" => 
-- sub_element <= PolyA(420);
        -- when "1001011000" => 
-- sub_element <= PolyA(419);
        -- when "1001011001" => 
-- sub_element <= PolyA(418);
        -- when "1001011010" => 
-- sub_element <= PolyA(417);
        -- when "1001011011" => 
-- sub_element <= PolyA(416);
        -- when "1001011100" => 
-- sub_element <= PolyA(415);
        -- when "1001011101" => 
-- sub_element <= PolyA(414);
        -- when "1001011110" => 
-- sub_element <= PolyA(413);
        -- when "1001011111" => 
-- sub_element <= PolyA(412);
        -- when "1001100000" => 
-- sub_element <= PolyA(411);
        -- when "1001100001" => 
-- sub_element <= PolyA(410);
        -- when "1001100010" => 
-- sub_element <= PolyA(409);
        -- when "1001100011" => 
-- sub_element <= PolyA(408);
        -- when "1001100100" => 
-- sub_element <= PolyA(407);
        -- when "1001100101" => 
-- sub_element <= PolyA(406);
        -- when "1001100110" => 
-- sub_element <= PolyA(405);
        -- when "1001100111" => 
-- sub_element <= PolyA(404);
        -- when "1001101000" => 
-- sub_element <= PolyA(403);
        -- when "1001101001" => 
-- sub_element <= PolyA(402);
        -- when "1001101010" => 
-- sub_element <= PolyA(401);
        -- when "1001101011" => 
-- sub_element <= PolyA(400);
        -- when "1001101100" => 
-- sub_element <= PolyA(399);
        -- when "1001101101" => 
-- sub_element <= PolyA(398);
        -- when "1001101110" => 
-- sub_element <= PolyA(397);
        -- when "1001101111" => 
-- sub_element <= PolyA(396);
        -- when "1001110000" => 
-- sub_element <= PolyA(395);
        -- when "1001110001" => 
-- sub_element <= PolyA(394);
        -- when "1001110010" => 
-- sub_element <= PolyA(393);
        -- when "1001110011" => 
-- sub_element <= PolyA(392);
        -- when "1001110100" => 
-- sub_element <= PolyA(391);
        -- when "1001110101" => 
-- sub_element <= PolyA(390);
        -- when "1001110110" => 
-- sub_element <= PolyA(389);
        -- when "1001110111" => 
-- sub_element <= PolyA(388);
        -- when "1001111000" => 
-- sub_element <= PolyA(387);
        -- when "1001111001" => 
-- sub_element <= PolyA(386);
        -- when "1001111010" => 
-- sub_element <= PolyA(385);
        -- when "1001111011" => 
-- sub_element <= PolyA(384);
        -- when "1001111100" => 
-- sub_element <= PolyA(383);
        -- when "1001111101" => 
-- sub_element <= PolyA(382);
        -- when "1001111110" => 
-- sub_element <= PolyA(381);
        -- when "1001111111" => 
-- sub_element <= PolyA(380);
        -- when "1010000000" => 
-- sub_element <= PolyA(379);
        -- when "1010000001" => 
-- sub_element <= PolyA(378);
        -- when "1010000010" => 
-- sub_element <= PolyA(377);
        -- when "1010000011" => 
-- sub_element <= PolyA(376);
        -- when "1010000100" => 
-- sub_element <= PolyA(375);
        -- when "1010000101" => 
-- sub_element <= PolyA(374);
        -- when "1010000110" => 
-- sub_element <= PolyA(373);
        -- when "1010000111" => 
-- sub_element <= PolyA(372);
        -- when "1010001000" => 
-- sub_element <= PolyA(371);
        -- when "1010001001" => 
-- sub_element <= PolyA(370);
        -- when "1010001010" => 
-- sub_element <= PolyA(369);
        -- when "1010001011" => 
-- sub_element <= PolyA(368);
        -- when "1010001100" => 
-- sub_element <= PolyA(367);
        -- when "1010001101" => 
-- sub_element <= PolyA(366);
        -- when "1010001110" => 
-- sub_element <= PolyA(365);
        -- when "1010001111" => 
-- sub_element <= PolyA(364);
        -- when "1010010000" => 
-- sub_element <= PolyA(363);
        -- when "1010010001" => 
-- sub_element <= PolyA(362);
        -- when "1010010010" => 
-- sub_element <= PolyA(361);
        -- when "1010010011" => 
-- sub_element <= PolyA(360);
        -- when "1010010100" => 
-- sub_element <= PolyA(359);
        -- when "1010010101" => 
-- sub_element <= PolyA(358);
        -- when "1010010110" => 
-- sub_element <= PolyA(357);
        -- when "1010010111" => 
-- sub_element <= PolyA(356);
        -- when "1010011000" => 
-- sub_element <= PolyA(355);
        -- when "1010011001" => 
-- sub_element <= PolyA(354);
        -- when "1010011010" => 
-- sub_element <= PolyA(353);
        -- when "1010011011" => 
-- sub_element <= PolyA(352);
        -- when "1010011100" => 
-- sub_element <= PolyA(351);
        -- when "1010011101" => 
-- sub_element <= PolyA(350);
        -- when "1010011110" => 
-- sub_element <= PolyA(349);
        -- when "1010011111" => 
-- sub_element <= PolyA(348);
        -- when "1010100000" => 
-- sub_element <= PolyA(347);
        -- when "1010100001" => 
-- sub_element <= PolyA(346);
        -- when "1010100010" => 
-- sub_element <= PolyA(345);
        -- when "1010100011" => 
-- sub_element <= PolyA(344);
        -- when "1010100100" => 
-- sub_element <= PolyA(343);
        -- when "1010100101" => 
-- sub_element <= PolyA(342);
        -- when "1010100110" => 
-- sub_element <= PolyA(341);
        -- when "1010100111" => 
-- sub_element <= PolyA(340);
        -- when "1010101000" => 
-- sub_element <= PolyA(339);
        -- when "1010101001" => 
-- sub_element <= PolyA(338);
        -- when "1010101010" => 
-- sub_element <= PolyA(337);
        -- when "1010101011" => 
-- sub_element <= PolyA(336);
        -- when "1010101100" => 
-- sub_element <= PolyA(335);
        -- when "1010101101" => 
-- sub_element <= PolyA(334);
        -- when "1010101110" => 
-- sub_element <= PolyA(333);
        -- when "1010101111" => 
-- sub_element <= PolyA(332);
        -- when "1010110000" => 
-- sub_element <= PolyA(331);
        -- when "1010110001" => 
-- sub_element <= PolyA(330);
        -- when "1010110010" => 
-- sub_element <= PolyA(329);
        -- when "1010110011" => 
-- sub_element <= PolyA(328);
        -- when "1010110100" => 
-- sub_element <= PolyA(327);
        -- when "1010110101" => 
-- sub_element <= PolyA(326);
        -- when "1010110110" => 
-- sub_element <= PolyA(325);
        -- when "1010110111" => 
-- sub_element <= PolyA(324);
        -- when "1010111000" => 
-- sub_element <= PolyA(323);
        -- when "1010111001" => 
-- sub_element <= PolyA(322);
        -- when "1010111010" => 
-- sub_element <= PolyA(321);
        -- when "1010111011" => 
-- sub_element <= PolyA(320);
        -- when "1010111100" => 
-- sub_element <= PolyA(319);
        -- when "1010111101" => 
-- sub_element <= PolyA(318);
        -- when "1010111110" => 
-- sub_element <= PolyA(317);
        -- when "1010111111" => 
-- sub_element <= PolyA(316);
        -- when "1011000000" => 
-- sub_element <= PolyA(315);
        -- when "1011000001" => 
-- sub_element <= PolyA(314);
        -- when "1011000010" => 
-- sub_element <= PolyA(313);
        -- when "1011000011" => 
-- sub_element <= PolyA(312);
        -- when "1011000100" => 
-- sub_element <= PolyA(311);
        -- when "1011000101" => 
-- sub_element <= PolyA(310);
        -- when "1011000110" => 
-- sub_element <= PolyA(309);
        -- when "1011000111" => 
-- sub_element <= PolyA(308);
        -- when "1011001000" => 
-- sub_element <= PolyA(307);
        -- when "1011001001" => 
-- sub_element <= PolyA(306);
        -- when "1011001010" => 
-- sub_element <= PolyA(305);
        -- when "1011001011" => 
-- sub_element <= PolyA(304);
        -- when "1011001100" => 
-- sub_element <= PolyA(303);
        -- when "1011001101" => 
-- sub_element <= PolyA(302);
        -- when "1011001110" => 
-- sub_element <= PolyA(301);
        -- when "1011001111" => 
-- sub_element <= PolyA(300);
        -- when "1011010000" => 
-- sub_element <= PolyA(299);
        -- when "1011010001" => 
-- sub_element <= PolyA(298);
        -- when "1011010010" => 
-- sub_element <= PolyA(297);
        -- when "1011010011" => 
-- sub_element <= PolyA(296);
        -- when "1011010100" => 
-- sub_element <= PolyA(295);
        -- when "1011010101" => 
-- sub_element <= PolyA(294);
        -- when "1011010110" => 
-- sub_element <= PolyA(293);
        -- when "1011010111" => 
-- sub_element <= PolyA(292);
        -- when "1011011000" => 
-- sub_element <= PolyA(291);
        -- when "1011011001" => 
-- sub_element <= PolyA(290);
        -- when "1011011010" => 
-- sub_element <= PolyA(289);
        -- when "1011011011" => 
-- sub_element <= PolyA(288);
        -- when "1011011100" => 
-- sub_element <= PolyA(287);
        -- when "1011011101" => 
-- sub_element <= PolyA(286);
        -- when "1011011110" => 
-- sub_element <= PolyA(285);
        -- when "1011011111" => 
-- sub_element <= PolyA(284);
        -- when "1011100000" => 
-- sub_element <= PolyA(283);
        -- when "1011100001" => 
-- sub_element <= PolyA(282);
        -- when "1011100010" => 
-- sub_element <= PolyA(281);
        -- when "1011100011" => 
-- sub_element <= PolyA(280);
        -- when "1011100100" => 
-- sub_element <= PolyA(279);
        -- when "1011100101" => 
-- sub_element <= PolyA(278);
        -- when "1011100110" => 
-- sub_element <= PolyA(277);
        -- when "1011100111" => 
-- sub_element <= PolyA(276);
        -- when "1011101000" => 
-- sub_element <= PolyA(275);
        -- when "1011101001" => 
-- sub_element <= PolyA(274);
        -- when "1011101010" => 
-- sub_element <= PolyA(273);
        -- when "1011101011" => 
-- sub_element <= PolyA(272);
        -- when "1011101100" => 
-- sub_element <= PolyA(271);
        -- when "1011101101" => 
-- sub_element <= PolyA(270);
        -- when "1011101110" => 
-- sub_element <= PolyA(269);
        -- when "1011101111" => 
-- sub_element <= PolyA(268);
        -- when "1011110000" => 
-- sub_element <= PolyA(267);
        -- when "1011110001" => 
-- sub_element <= PolyA(266);
        -- when "1011110010" => 
-- sub_element <= PolyA(265);
        -- when "1011110011" => 
-- sub_element <= PolyA(264);
        -- when "1011110100" => 
-- sub_element <= PolyA(263);
        -- when "1011110101" => 
-- sub_element <= PolyA(262);
        -- when "1011110110" => 
-- sub_element <= PolyA(261);
        -- when "1011110111" => 
-- sub_element <= PolyA(260);
        -- when "1011111000" => 
-- sub_element <= PolyA(259);
        -- when "1011111001" => 
-- sub_element <= PolyA(258);
        -- when "1011111010" => 
-- sub_element <= PolyA(257);
        -- when "1011111011" => 
-- sub_element <= PolyA(256);
        -- when "1011111100" => 
-- sub_element <= PolyA(255);
        -- when "1011111101" => 
-- sub_element <= PolyA(254);
        -- when "1011111110" => 
-- sub_element <= PolyA(253);
        -- when "1011111111" => 
-- sub_element <= PolyA(252);
        -- when "1100000000" => 
-- sub_element <= PolyA(251);
        -- when "1100000001" => 
-- sub_element <= PolyA(250);
        -- when "1100000010" => 
-- sub_element <= PolyA(249);
        -- when "1100000011" => 
-- sub_element <= PolyA(248);
        -- when "1100000100" => 
-- sub_element <= PolyA(247);
        -- when "1100000101" => 
-- sub_element <= PolyA(246);
        -- when "1100000110" => 
-- sub_element <= PolyA(245);
        -- when "1100000111" => 
-- sub_element <= PolyA(244);
        -- when "1100001000" => 
-- sub_element <= PolyA(243);
        -- when "1100001001" => 
-- sub_element <= PolyA(242);
        -- when "1100001010" => 
-- sub_element <= PolyA(241);
        -- when "1100001011" => 
-- sub_element <= PolyA(240);
        -- when "1100001100" => 
-- sub_element <= PolyA(239);
        -- when "1100001101" => 
-- sub_element <= PolyA(238);
        -- when "1100001110" => 
-- sub_element <= PolyA(237);
        -- when "1100001111" => 
-- sub_element <= PolyA(236);
        -- when "1100010000" => 
-- sub_element <= PolyA(235);
        -- when "1100010001" => 
-- sub_element <= PolyA(234);
        -- when "1100010010" => 
-- sub_element <= PolyA(233);
        -- when "1100010011" => 
-- sub_element <= PolyA(232);
        -- when "1100010100" => 
-- sub_element <= PolyA(231);
        -- when "1100010101" => 
-- sub_element <= PolyA(230);
        -- when "1100010110" => 
-- sub_element <= PolyA(229);
        -- when "1100010111" => 
-- sub_element <= PolyA(228);
        -- when "1100011000" => 
-- sub_element <= PolyA(227);
        -- when "1100011001" => 
-- sub_element <= PolyA(226);
        -- when "1100011010" => 
-- sub_element <= PolyA(225);
        -- when "1100011011" => 
-- sub_element <= PolyA(224);
        -- when "1100011100" => 
-- sub_element <= PolyA(223);
        -- when "1100011101" => 
-- sub_element <= PolyA(222);
        -- when "1100011110" => 
-- sub_element <= PolyA(221);
        -- when "1100011111" => 
-- sub_element <= PolyA(220);
        -- when "1100100000" => 
-- sub_element <= PolyA(219);
        -- when "1100100001" => 
-- sub_element <= PolyA(218);
        -- when "1100100010" => 
-- sub_element <= PolyA(217);
        -- when "1100100011" => 
-- sub_element <= PolyA(216);
        -- when "1100100100" => 
-- sub_element <= PolyA(215);
        -- when "1100100101" => 
-- sub_element <= PolyA(214);
        -- when "1100100110" => 
-- sub_element <= PolyA(213);
        -- when "1100100111" => 
-- sub_element <= PolyA(212);
        -- when "1100101000" => 
-- sub_element <= PolyA(211);
        -- when "1100101001" => 
-- sub_element <= PolyA(210);
        -- when "1100101010" => 
-- sub_element <= PolyA(209);
        -- when "1100101011" => 
-- sub_element <= PolyA(208);
        -- when "1100101100" => 
-- sub_element <= PolyA(207);
        -- when "1100101101" => 
-- sub_element <= PolyA(206);
        -- when "1100101110" => 
-- sub_element <= PolyA(205);
        -- when "1100101111" => 
-- sub_element <= PolyA(204);
        -- when "1100110000" => 
-- sub_element <= PolyA(203);
        -- when "1100110001" => 
-- sub_element <= PolyA(202);
        -- when "1100110010" => 
-- sub_element <= PolyA(201);
        -- when "1100110011" => 
-- sub_element <= PolyA(200);
        -- when "1100110100" => 
-- sub_element <= PolyA(199);
        -- when "1100110101" => 
-- sub_element <= PolyA(198);
        -- when "1100110110" => 
-- sub_element <= PolyA(197);
        -- when "1100110111" => 
-- sub_element <= PolyA(196);
        -- when "1100111000" => 
-- sub_element <= PolyA(195);
        -- when "1100111001" => 
-- sub_element <= PolyA(194);
        -- when "1100111010" => 
-- sub_element <= PolyA(193);
        -- when "1100111011" => 
-- sub_element <= PolyA(192);
        -- when "1100111100" => 
-- sub_element <= PolyA(191);
        -- when "1100111101" => 
-- sub_element <= PolyA(190);
        -- when "1100111110" => 
-- sub_element <= PolyA(189);
        -- when "1100111111" => 
-- sub_element <= PolyA(188);
        -- when "1101000000" => 
-- sub_element <= PolyA(187);
        -- when "1101000001" => 
-- sub_element <= PolyA(186);
        -- when "1101000010" => 
-- sub_element <= PolyA(185);
        -- when "1101000011" => 
-- sub_element <= PolyA(184);
        -- when "1101000100" => 
-- sub_element <= PolyA(183);
        -- when "1101000101" => 
-- sub_element <= PolyA(182);
        -- when "1101000110" => 
-- sub_element <= PolyA(181);
        -- when "1101000111" => 
-- sub_element <= PolyA(180);
        -- when "1101001000" => 
-- sub_element <= PolyA(179);
        -- when "1101001001" => 
-- sub_element <= PolyA(178);
        -- when "1101001010" => 
-- sub_element <= PolyA(177);
        -- when "1101001011" => 
-- sub_element <= PolyA(176);
        -- when "1101001100" => 
-- sub_element <= PolyA(175);
        -- when "1101001101" => 
-- sub_element <= PolyA(174);
        -- when "1101001110" => 
-- sub_element <= PolyA(173);
        -- when "1101001111" => 
-- sub_element <= PolyA(172);
        -- when "1101010000" => 
-- sub_element <= PolyA(171);
        -- when "1101010001" => 
-- sub_element <= PolyA(170);
        -- when "1101010010" => 
-- sub_element <= PolyA(169);
        -- when "1101010011" => 
-- sub_element <= PolyA(168);
        -- when "1101010100" => 
-- sub_element <= PolyA(167);
        -- when "1101010101" => 
-- sub_element <= PolyA(166);
        -- when "1101010110" => 
-- sub_element <= PolyA(165);
        -- when "1101010111" => 
-- sub_element <= PolyA(164);
        -- when "1101011000" => 
-- sub_element <= PolyA(163);
        -- when "1101011001" => 
-- sub_element <= PolyA(162);
        -- when "1101011010" => 
-- sub_element <= PolyA(161);
        -- when "1101011011" => 
-- sub_element <= PolyA(160);
        -- when "1101011100" => 
-- sub_element <= PolyA(159);
        -- when "1101011101" => 
-- sub_element <= PolyA(158);
        -- when "1101011110" => 
-- sub_element <= PolyA(157);
        -- when "1101011111" => 
-- sub_element <= PolyA(156);
        -- when "1101100000" => 
-- sub_element <= PolyA(155);
        -- when "1101100001" => 
-- sub_element <= PolyA(154);
        -- when "1101100010" => 
-- sub_element <= PolyA(153);
        -- when "1101100011" => 
-- sub_element <= PolyA(152);
        -- when "1101100100" => 
-- sub_element <= PolyA(151);
        -- when "1101100101" => 
-- sub_element <= PolyA(150);
        -- when "1101100110" => 
-- sub_element <= PolyA(149);
        -- when "1101100111" => 
-- sub_element <= PolyA(148);
        -- when "1101101000" => 
-- sub_element <= PolyA(147);
        -- when "1101101001" => 
-- sub_element <= PolyA(146);
        -- when "1101101010" => 
-- sub_element <= PolyA(145);
        -- when "1101101011" => 
-- sub_element <= PolyA(144);
        -- when "1101101100" => 
-- sub_element <= PolyA(143);
        -- when "1101101101" => 
-- sub_element <= PolyA(142);
        -- when "1101101110" => 
-- sub_element <= PolyA(141);
        -- when "1101101111" => 
-- sub_element <= PolyA(140);
        -- when "1101110000" => 
-- sub_element <= PolyA(139);
        -- when "1101110001" => 
-- sub_element <= PolyA(138);
        -- when "1101110010" => 
-- sub_element <= PolyA(137);
        -- when "1101110011" => 
-- sub_element <= PolyA(136);
        -- when "1101110100" => 
-- sub_element <= PolyA(135);
        -- when "1101110101" => 
-- sub_element <= PolyA(134);
        -- when "1101110110" => 
-- sub_element <= PolyA(133);
        -- when "1101110111" => 
-- sub_element <= PolyA(132);
        -- when "1101111000" => 
-- sub_element <= PolyA(131);
        -- when "1101111001" => 
-- sub_element <= PolyA(130);
        -- when "1101111010" => 
-- sub_element <= PolyA(129);
        -- when "1101111011" => 
-- sub_element <= PolyA(128);
        -- when "1101111100" => 
-- sub_element <= PolyA(127);
        -- when "1101111101" => 
-- sub_element <= PolyA(126);
        -- when "1101111110" => 
-- sub_element <= PolyA(125);
        -- when "1101111111" => 
-- sub_element <= PolyA(124);
        -- when "1110000000" => 
-- sub_element <= PolyA(123);
        -- when "1110000001" => 
-- sub_element <= PolyA(122);
        -- when "1110000010" => 
-- sub_element <= PolyA(121);
        -- when "1110000011" => 
-- sub_element <= PolyA(120);
        -- when "1110000100" => 
-- sub_element <= PolyA(119);
        -- when "1110000101" => 
-- sub_element <= PolyA(118);
        -- when "1110000110" => 
-- sub_element <= PolyA(117);
        -- when "1110000111" => 
-- sub_element <= PolyA(116);
        -- when "1110001000" => 
-- sub_element <= PolyA(115);
        -- when "1110001001" => 
-- sub_element <= PolyA(114);
        -- when "1110001010" => 
-- sub_element <= PolyA(113);
        -- when "1110001011" => 
-- sub_element <= PolyA(112);
        -- when "1110001100" => 
-- sub_element <= PolyA(111);
        -- when "1110001101" => 
-- sub_element <= PolyA(110);
        -- when "1110001110" => 
-- sub_element <= PolyA(109);
        -- when "1110001111" => 
-- sub_element <= PolyA(108);
        -- when "1110010000" => 
-- sub_element <= PolyA(107);
        -- when "1110010001" => 
-- sub_element <= PolyA(106);
        -- when "1110010010" => 
-- sub_element <= PolyA(105);
        -- when "1110010011" => 
-- sub_element <= PolyA(104);
        -- when "1110010100" => 
-- sub_element <= PolyA(103);
        -- when "1110010101" => 
-- sub_element <= PolyA(102);
        -- when "1110010110" => 
-- sub_element <= PolyA(101);
        -- when "1110010111" => 
-- sub_element <= PolyA(100);
        -- when "1110011000" => 
-- sub_element <= PolyA(99);
        -- when "1110011001" => 
-- sub_element <= PolyA(98);
        -- when "1110011010" => 
-- sub_element <= PolyA(97);
        -- when "1110011011" => 
-- sub_element <= PolyA(96);
        -- when "1110011100" => 
-- sub_element <= PolyA(95);
        -- when "1110011101" => 
-- sub_element <= PolyA(94);
        -- when "1110011110" => 
-- sub_element <= PolyA(93);
        -- when "1110011111" => 
-- sub_element <= PolyA(92);
        -- when "1110100000" => 
-- sub_element <= PolyA(91);
        -- when "1110100001" => 
-- sub_element <= PolyA(90);
        -- when "1110100010" => 
-- sub_element <= PolyA(89);
        -- when "1110100011" => 
-- sub_element <= PolyA(88);
        -- when "1110100100" => 
-- sub_element <= PolyA(87);
        -- when "1110100101" => 
-- sub_element <= PolyA(86);
        -- when "1110100110" => 
-- sub_element <= PolyA(85);
        -- when "1110100111" => 
-- sub_element <= PolyA(84);
        -- when "1110101000" => 
-- sub_element <= PolyA(83);
        -- when "1110101001" => 
-- sub_element <= PolyA(82);
        -- when "1110101010" => 
-- sub_element <= PolyA(81);
        -- when "1110101011" => 
-- sub_element <= PolyA(80);
        -- when "1110101100" => 
-- sub_element <= PolyA(79);
        -- when "1110101101" => 
-- sub_element <= PolyA(78);
        -- when "1110101110" => 
-- sub_element <= PolyA(77);
        -- when "1110101111" => 
-- sub_element <= PolyA(76);
        -- when "1110110000" => 
-- sub_element <= PolyA(75);
        -- when "1110110001" => 
-- sub_element <= PolyA(74);
        -- when "1110110010" => 
-- sub_element <= PolyA(73);
        -- when "1110110011" => 
-- sub_element <= PolyA(72);
        -- when "1110110100" => 
-- sub_element <= PolyA(71);
        -- when "1110110101" => 
-- sub_element <= PolyA(70);
        -- when "1110110110" => 
-- sub_element <= PolyA(69);
        -- when "1110110111" => 
-- sub_element <= PolyA(68);
        -- when "1110111000" => 
-- sub_element <= PolyA(67);
        -- when "1110111001" => 
-- sub_element <= PolyA(66);
        -- when "1110111010" => 
-- sub_element <= PolyA(65);
        -- when "1110111011" => 
-- sub_element <= PolyA(64);
        -- when "1110111100" => 
-- sub_element <= PolyA(63);
        -- when "1110111101" => 
-- sub_element <= PolyA(62);
        -- when "1110111110" => 
-- sub_element <= PolyA(61);
        -- when "1110111111" => 
-- sub_element <= PolyA(60);
        -- when "1111000000" => 
-- sub_element <= PolyA(59);
        -- when "1111000001" => 
-- sub_element <= PolyA(58);
        -- when "1111000010" => 
-- sub_element <= PolyA(57);
        -- when "1111000011" => 
-- sub_element <= PolyA(56);
        -- when "1111000100" => 
-- sub_element <= PolyA(55);
        -- when "1111000101" => 
-- sub_element <= PolyA(54);
        -- when "1111000110" => 
-- sub_element <= PolyA(53);
        -- when "1111000111" => 
-- sub_element <= PolyA(52);
        -- when "1111001000" => 
-- sub_element <= PolyA(51);
        -- when "1111001001" => 
-- sub_element <= PolyA(50);
        -- when "1111001010" => 
-- sub_element <= PolyA(49);
        -- when "1111001011" => 
-- sub_element <= PolyA(48);
        -- when "1111001100" => 
-- sub_element <= PolyA(47);
        -- when "1111001101" => 
-- sub_element <= PolyA(46);
        -- when "1111001110" => 
-- sub_element <= PolyA(45);
        -- when "1111001111" => 
-- sub_element <= PolyA(44);
        -- when "1111010000" => 
-- sub_element <= PolyA(43);
        -- when "1111010001" => 
-- sub_element <= PolyA(42);
        -- when "1111010010" => 
-- sub_element <= PolyA(41);
        -- when "1111010011" => 
-- sub_element <= PolyA(40);
        -- when "1111010100" => 
-- sub_element <= PolyA(39);
        -- when "1111010101" => 
-- sub_element <= PolyA(38);
        -- when "1111010110" => 
-- sub_element <= PolyA(37);
        -- when "1111010111" => 
-- sub_element <= PolyA(36);
        -- when "1111011000" => 
-- sub_element <= PolyA(35);
        -- when "1111011001" => 
-- sub_element <= PolyA(34);
        -- when "1111011010" => 
-- sub_element <= PolyA(33);
        -- when "1111011011" => 
-- sub_element <= PolyA(32);
        -- when "1111011100" => 
-- sub_element <= PolyA(31);
        -- when "1111011101" => 
-- sub_element <= PolyA(30);
        -- when "1111011110" => 
-- sub_element <= PolyA(29);
        -- when "1111011111" => 
-- sub_element <= PolyA(28);
        -- when "1111100000" => 
-- sub_element <= PolyA(27);
        -- when "1111100001" => 
-- sub_element <= PolyA(26);
        -- when "1111100010" => 
-- sub_element <= PolyA(25);
        -- when "1111100011" => 
-- sub_element <= PolyA(24);
        -- when "1111100100" => 
-- sub_element <= PolyA(23);
        -- when "1111100101" => 
-- sub_element <= PolyA(22);
        -- when "1111100110" => 
-- sub_element <= PolyA(21);
        -- when "1111100111" => 
-- sub_element <= PolyA(20);
        -- when "1111101000" => 
-- sub_element <= PolyA(19);
        -- when "1111101001" => 
-- sub_element <= PolyA(18);
        -- when "1111101010" => 
-- sub_element <= PolyA(17);
        -- when "1111101011" => 
-- sub_element <= PolyA(16);
        -- when "1111101100" => 
-- sub_element <= PolyA(15);
        -- when "1111101101" => 
-- sub_element <= PolyA(14);
        -- when "1111101110" => 
-- sub_element <= PolyA(13);
        -- when "1111101111" => 
-- sub_element <= PolyA(12);
        -- when "1111110000" => 
-- sub_element <= PolyA(11);
        -- when "1111110001" => 
-- sub_element <= PolyA(10);
        -- when "1111110010" => 
-- sub_element <= PolyA(9);
        -- when "1111110011" => 
-- sub_element <= PolyA(8);
        -- when "1111110100" => 
-- sub_element <= PolyA(7);
        -- when "1111110101" => 
-- sub_element <= PolyA(6);
        -- when "1111110110" => 
-- sub_element <= PolyA(5);
        -- when "1111110111" => 
-- sub_element <= PolyA(4);
        -- when "1111111000" => 
-- sub_element <= PolyA(3);
        -- when "1111111001" => 
-- sub_element <= PolyA(2);
        -- when "1111111010" => 
-- sub_element <= PolyA(1);
        -- when "1111111011" => 
-- sub_element <= PolyA(0);
         -- when others =>
             -- sub_element <= (others => '0');
     -- end case;
 -- end if;
-- end process;
----==========   OutPUT Pointer  ================
-- process(clk)
-- begin
 -- if clk'event and clk = '1' then
     -- case input_pointer is

        -- when "0000000010" => 
-- LongRes(1018) <= sub_result;
        -- when "0000000011" => 
-- LongRes(1017) <= sub_result;
        -- when "0000000100" => 
-- LongRes(1016) <= sub_result;
        -- when "0000000101" => 
-- LongRes(1015) <= sub_result;
        -- when "0000000110" => 
-- LongRes(1014) <= sub_result;
        -- when "0000000111" => 
-- LongRes(1013) <= sub_result;
        -- when "0000001000" => 
-- LongRes(1012) <= sub_result;
        -- when "0000001001" => 
-- LongRes(1011) <= sub_result;
        -- when "0000001010" => 
-- LongRes(1010) <= sub_result;
        -- when "0000001011" => 
-- LongRes(1009) <= sub_result;
        -- when "0000001100" => 
-- LongRes(1008) <= sub_result;
        -- when "0000001101" => 
-- LongRes(1007) <= sub_result;
        -- when "0000001110" => 
-- LongRes(1006) <= sub_result;
        -- when "0000001111" => 
-- LongRes(1005) <= sub_result;
        -- when "0000010000" => 
-- LongRes(1004) <= sub_result;
        -- when "0000010001" => 
-- LongRes(1003) <= sub_result;
        -- when "0000010010" => 
-- LongRes(1002) <= sub_result;
        -- when "0000010011" => 
-- LongRes(1001) <= sub_result;
        -- when "0000010100" => 
-- LongRes(1000) <= sub_result;
        -- when "0000010101" => 
-- LongRes(999) <= sub_result;
        -- when "0000010110" => 
-- LongRes(998) <= sub_result;
        -- when "0000010111" => 
-- LongRes(997) <= sub_result;
        -- when "0000011000" => 
-- LongRes(996) <= sub_result;
        -- when "0000011001" => 
-- LongRes(995) <= sub_result;
        -- when "0000011010" => 
-- LongRes(994) <= sub_result;
        -- when "0000011011" => 
-- LongRes(993) <= sub_result;
        -- when "0000011100" => 
-- LongRes(992) <= sub_result;
        -- when "0000011101" => 
-- LongRes(991) <= sub_result;
        -- when "0000011110" => 
-- LongRes(990) <= sub_result;
        -- when "0000011111" => 
-- LongRes(989) <= sub_result;
        -- when "0000100000" => 
-- LongRes(988) <= sub_result;
        -- when "0000100001" => 
-- LongRes(987) <= sub_result;
        -- when "0000100010" => 
-- LongRes(986) <= sub_result;
        -- when "0000100011" => 
-- LongRes(985) <= sub_result;
        -- when "0000100100" => 
-- LongRes(984) <= sub_result;
        -- when "0000100101" => 
-- LongRes(983) <= sub_result;
        -- when "0000100110" => 
-- LongRes(982) <= sub_result;
        -- when "0000100111" => 
-- LongRes(981) <= sub_result;
        -- when "0000101000" => 
-- LongRes(980) <= sub_result;
        -- when "0000101001" => 
-- LongRes(979) <= sub_result;
        -- when "0000101010" => 
-- LongRes(978) <= sub_result;
        -- when "0000101011" => 
-- LongRes(977) <= sub_result;
        -- when "0000101100" => 
-- LongRes(976) <= sub_result;
        -- when "0000101101" => 
-- LongRes(975) <= sub_result;
        -- when "0000101110" => 
-- LongRes(974) <= sub_result;
        -- when "0000101111" => 
-- LongRes(973) <= sub_result;
        -- when "0000110000" => 
-- LongRes(972) <= sub_result;
        -- when "0000110001" => 
-- LongRes(971) <= sub_result;
        -- when "0000110010" => 
-- LongRes(970) <= sub_result;
        -- when "0000110011" => 
-- LongRes(969) <= sub_result;
        -- when "0000110100" => 
-- LongRes(968) <= sub_result;
        -- when "0000110101" => 
-- LongRes(967) <= sub_result;
        -- when "0000110110" => 
-- LongRes(966) <= sub_result;
        -- when "0000110111" => 
-- LongRes(965) <= sub_result;
        -- when "0000111000" => 
-- LongRes(964) <= sub_result;
        -- when "0000111001" => 
-- LongRes(963) <= sub_result;
        -- when "0000111010" => 
-- LongRes(962) <= sub_result;
        -- when "0000111011" => 
-- LongRes(961) <= sub_result;
        -- when "0000111100" => 
-- LongRes(960) <= sub_result;
        -- when "0000111101" => 
-- LongRes(959) <= sub_result;
        -- when "0000111110" => 
-- LongRes(958) <= sub_result;
        -- when "0000111111" => 
-- LongRes(957) <= sub_result;
        -- when "0001000000" => 
-- LongRes(956) <= sub_result;
        -- when "0001000001" => 
-- LongRes(955) <= sub_result;
        -- when "0001000010" => 
-- LongRes(954) <= sub_result;
        -- when "0001000011" => 
-- LongRes(953) <= sub_result;
        -- when "0001000100" => 
-- LongRes(952) <= sub_result;
        -- when "0001000101" => 
-- LongRes(951) <= sub_result;
        -- when "0001000110" => 
-- LongRes(950) <= sub_result;
        -- when "0001000111" => 
-- LongRes(949) <= sub_result;
        -- when "0001001000" => 
-- LongRes(948) <= sub_result;
        -- when "0001001001" => 
-- LongRes(947) <= sub_result;
        -- when "0001001010" => 
-- LongRes(946) <= sub_result;
        -- when "0001001011" => 
-- LongRes(945) <= sub_result;
        -- when "0001001100" => 
-- LongRes(944) <= sub_result;
        -- when "0001001101" => 
-- LongRes(943) <= sub_result;
        -- when "0001001110" => 
-- LongRes(942) <= sub_result;
        -- when "0001001111" => 
-- LongRes(941) <= sub_result;
        -- when "0001010000" => 
-- LongRes(940) <= sub_result;
        -- when "0001010001" => 
-- LongRes(939) <= sub_result;
        -- when "0001010010" => 
-- LongRes(938) <= sub_result;
        -- when "0001010011" => 
-- LongRes(937) <= sub_result;
        -- when "0001010100" => 
-- LongRes(936) <= sub_result;
        -- when "0001010101" => 
-- LongRes(935) <= sub_result;
        -- when "0001010110" => 
-- LongRes(934) <= sub_result;
        -- when "0001010111" => 
-- LongRes(933) <= sub_result;
        -- when "0001011000" => 
-- LongRes(932) <= sub_result;
        -- when "0001011001" => 
-- LongRes(931) <= sub_result;
        -- when "0001011010" => 
-- LongRes(930) <= sub_result;
        -- when "0001011011" => 
-- LongRes(929) <= sub_result;
        -- when "0001011100" => 
-- LongRes(928) <= sub_result;
        -- when "0001011101" => 
-- LongRes(927) <= sub_result;
        -- when "0001011110" => 
-- LongRes(926) <= sub_result;
        -- when "0001011111" => 
-- LongRes(925) <= sub_result;
        -- when "0001100000" => 
-- LongRes(924) <= sub_result;
        -- when "0001100001" => 
-- LongRes(923) <= sub_result;
        -- when "0001100010" => 
-- LongRes(922) <= sub_result;
        -- when "0001100011" => 
-- LongRes(921) <= sub_result;
        -- when "0001100100" => 
-- LongRes(920) <= sub_result;
        -- when "0001100101" => 
-- LongRes(919) <= sub_result;
        -- when "0001100110" => 
-- LongRes(918) <= sub_result;
        -- when "0001100111" => 
-- LongRes(917) <= sub_result;
        -- when "0001101000" => 
-- LongRes(916) <= sub_result;
        -- when "0001101001" => 
-- LongRes(915) <= sub_result;
        -- when "0001101010" => 
-- LongRes(914) <= sub_result;
        -- when "0001101011" => 
-- LongRes(913) <= sub_result;
        -- when "0001101100" => 
-- LongRes(912) <= sub_result;
        -- when "0001101101" => 
-- LongRes(911) <= sub_result;
        -- when "0001101110" => 
-- LongRes(910) <= sub_result;
        -- when "0001101111" => 
-- LongRes(909) <= sub_result;
        -- when "0001110000" => 
-- LongRes(908) <= sub_result;
        -- when "0001110001" => 
-- LongRes(907) <= sub_result;
        -- when "0001110010" => 
-- LongRes(906) <= sub_result;
        -- when "0001110011" => 
-- LongRes(905) <= sub_result;
        -- when "0001110100" => 
-- LongRes(904) <= sub_result;
        -- when "0001110101" => 
-- LongRes(903) <= sub_result;
        -- when "0001110110" => 
-- LongRes(902) <= sub_result;
        -- when "0001110111" => 
-- LongRes(901) <= sub_result;
        -- when "0001111000" => 
-- LongRes(900) <= sub_result;
        -- when "0001111001" => 
-- LongRes(899) <= sub_result;
        -- when "0001111010" => 
-- LongRes(898) <= sub_result;
        -- when "0001111011" => 
-- LongRes(897) <= sub_result;
        -- when "0001111100" => 
-- LongRes(896) <= sub_result;
        -- when "0001111101" => 
-- LongRes(895) <= sub_result;
        -- when "0001111110" => 
-- LongRes(894) <= sub_result;
        -- when "0001111111" => 
-- LongRes(893) <= sub_result;
        -- when "0010000000" => 
-- LongRes(892) <= sub_result;
        -- when "0010000001" => 
-- LongRes(891) <= sub_result;
        -- when "0010000010" => 
-- LongRes(890) <= sub_result;
        -- when "0010000011" => 
-- LongRes(889) <= sub_result;
        -- when "0010000100" => 
-- LongRes(888) <= sub_result;
        -- when "0010000101" => 
-- LongRes(887) <= sub_result;
        -- when "0010000110" => 
-- LongRes(886) <= sub_result;
        -- when "0010000111" => 
-- LongRes(885) <= sub_result;
        -- when "0010001000" => 
-- LongRes(884) <= sub_result;
        -- when "0010001001" => 
-- LongRes(883) <= sub_result;
        -- when "0010001010" => 
-- LongRes(882) <= sub_result;
        -- when "0010001011" => 
-- LongRes(881) <= sub_result;
        -- when "0010001100" => 
-- LongRes(880) <= sub_result;
        -- when "0010001101" => 
-- LongRes(879) <= sub_result;
        -- when "0010001110" => 
-- LongRes(878) <= sub_result;
        -- when "0010001111" => 
-- LongRes(877) <= sub_result;
        -- when "0010010000" => 
-- LongRes(876) <= sub_result;
        -- when "0010010001" => 
-- LongRes(875) <= sub_result;
        -- when "0010010010" => 
-- LongRes(874) <= sub_result;
        -- when "0010010011" => 
-- LongRes(873) <= sub_result;
        -- when "0010010100" => 
-- LongRes(872) <= sub_result;
        -- when "0010010101" => 
-- LongRes(871) <= sub_result;
        -- when "0010010110" => 
-- LongRes(870) <= sub_result;
        -- when "0010010111" => 
-- LongRes(869) <= sub_result;
        -- when "0010011000" => 
-- LongRes(868) <= sub_result;
        -- when "0010011001" => 
-- LongRes(867) <= sub_result;
        -- when "0010011010" => 
-- LongRes(866) <= sub_result;
        -- when "0010011011" => 
-- LongRes(865) <= sub_result;
        -- when "0010011100" => 
-- LongRes(864) <= sub_result;
        -- when "0010011101" => 
-- LongRes(863) <= sub_result;
        -- when "0010011110" => 
-- LongRes(862) <= sub_result;
        -- when "0010011111" => 
-- LongRes(861) <= sub_result;
        -- when "0010100000" => 
-- LongRes(860) <= sub_result;
        -- when "0010100001" => 
-- LongRes(859) <= sub_result;
        -- when "0010100010" => 
-- LongRes(858) <= sub_result;
        -- when "0010100011" => 
-- LongRes(857) <= sub_result;
        -- when "0010100100" => 
-- LongRes(856) <= sub_result;
        -- when "0010100101" => 
-- LongRes(855) <= sub_result;
        -- when "0010100110" => 
-- LongRes(854) <= sub_result;
        -- when "0010100111" => 
-- LongRes(853) <= sub_result;
        -- when "0010101000" => 
-- LongRes(852) <= sub_result;
        -- when "0010101001" => 
-- LongRes(851) <= sub_result;
        -- when "0010101010" => 
-- LongRes(850) <= sub_result;
        -- when "0010101011" => 
-- LongRes(849) <= sub_result;
        -- when "0010101100" => 
-- LongRes(848) <= sub_result;
        -- when "0010101101" => 
-- LongRes(847) <= sub_result;
        -- when "0010101110" => 
-- LongRes(846) <= sub_result;
        -- when "0010101111" => 
-- LongRes(845) <= sub_result;
        -- when "0010110000" => 
-- LongRes(844) <= sub_result;
        -- when "0010110001" => 
-- LongRes(843) <= sub_result;
        -- when "0010110010" => 
-- LongRes(842) <= sub_result;
        -- when "0010110011" => 
-- LongRes(841) <= sub_result;
        -- when "0010110100" => 
-- LongRes(840) <= sub_result;
        -- when "0010110101" => 
-- LongRes(839) <= sub_result;
        -- when "0010110110" => 
-- LongRes(838) <= sub_result;
        -- when "0010110111" => 
-- LongRes(837) <= sub_result;
        -- when "0010111000" => 
-- LongRes(836) <= sub_result;
        -- when "0010111001" => 
-- LongRes(835) <= sub_result;
        -- when "0010111010" => 
-- LongRes(834) <= sub_result;
        -- when "0010111011" => 
-- LongRes(833) <= sub_result;
        -- when "0010111100" => 
-- LongRes(832) <= sub_result;
        -- when "0010111101" => 
-- LongRes(831) <= sub_result;
        -- when "0010111110" => 
-- LongRes(830) <= sub_result;
        -- when "0010111111" => 
-- LongRes(829) <= sub_result;
        -- when "0011000000" => 
-- LongRes(828) <= sub_result;
        -- when "0011000001" => 
-- LongRes(827) <= sub_result;
        -- when "0011000010" => 
-- LongRes(826) <= sub_result;
        -- when "0011000011" => 
-- LongRes(825) <= sub_result;
        -- when "0011000100" => 
-- LongRes(824) <= sub_result;
        -- when "0011000101" => 
-- LongRes(823) <= sub_result;
        -- when "0011000110" => 
-- LongRes(822) <= sub_result;
        -- when "0011000111" => 
-- LongRes(821) <= sub_result;
        -- when "0011001000" => 
-- LongRes(820) <= sub_result;
        -- when "0011001001" => 
-- LongRes(819) <= sub_result;
        -- when "0011001010" => 
-- LongRes(818) <= sub_result;
        -- when "0011001011" => 
-- LongRes(817) <= sub_result;
        -- when "0011001100" => 
-- LongRes(816) <= sub_result;
        -- when "0011001101" => 
-- LongRes(815) <= sub_result;
        -- when "0011001110" => 
-- LongRes(814) <= sub_result;
        -- when "0011001111" => 
-- LongRes(813) <= sub_result;
        -- when "0011010000" => 
-- LongRes(812) <= sub_result;
        -- when "0011010001" => 
-- LongRes(811) <= sub_result;
        -- when "0011010010" => 
-- LongRes(810) <= sub_result;
        -- when "0011010011" => 
-- LongRes(809) <= sub_result;
        -- when "0011010100" => 
-- LongRes(808) <= sub_result;
        -- when "0011010101" => 
-- LongRes(807) <= sub_result;
        -- when "0011010110" => 
-- LongRes(806) <= sub_result;
        -- when "0011010111" => 
-- LongRes(805) <= sub_result;
        -- when "0011011000" => 
-- LongRes(804) <= sub_result;
        -- when "0011011001" => 
-- LongRes(803) <= sub_result;
        -- when "0011011010" => 
-- LongRes(802) <= sub_result;
        -- when "0011011011" => 
-- LongRes(801) <= sub_result;
        -- when "0011011100" => 
-- LongRes(800) <= sub_result;
        -- when "0011011101" => 
-- LongRes(799) <= sub_result;
        -- when "0011011110" => 
-- LongRes(798) <= sub_result;
        -- when "0011011111" => 
-- LongRes(797) <= sub_result;
        -- when "0011100000" => 
-- LongRes(796) <= sub_result;
        -- when "0011100001" => 
-- LongRes(795) <= sub_result;
        -- when "0011100010" => 
-- LongRes(794) <= sub_result;
        -- when "0011100011" => 
-- LongRes(793) <= sub_result;
        -- when "0011100100" => 
-- LongRes(792) <= sub_result;
        -- when "0011100101" => 
-- LongRes(791) <= sub_result;
        -- when "0011100110" => 
-- LongRes(790) <= sub_result;
        -- when "0011100111" => 
-- LongRes(789) <= sub_result;
        -- when "0011101000" => 
-- LongRes(788) <= sub_result;
        -- when "0011101001" => 
-- LongRes(787) <= sub_result;
        -- when "0011101010" => 
-- LongRes(786) <= sub_result;
        -- when "0011101011" => 
-- LongRes(785) <= sub_result;
        -- when "0011101100" => 
-- LongRes(784) <= sub_result;
        -- when "0011101101" => 
-- LongRes(783) <= sub_result;
        -- when "0011101110" => 
-- LongRes(782) <= sub_result;
        -- when "0011101111" => 
-- LongRes(781) <= sub_result;
        -- when "0011110000" => 
-- LongRes(780) <= sub_result;
        -- when "0011110001" => 
-- LongRes(779) <= sub_result;
        -- when "0011110010" => 
-- LongRes(778) <= sub_result;
        -- when "0011110011" => 
-- LongRes(777) <= sub_result;
        -- when "0011110100" => 
-- LongRes(776) <= sub_result;
        -- when "0011110101" => 
-- LongRes(775) <= sub_result;
        -- when "0011110110" => 
-- LongRes(774) <= sub_result;
        -- when "0011110111" => 
-- LongRes(773) <= sub_result;
        -- when "0011111000" => 
-- LongRes(772) <= sub_result;
        -- when "0011111001" => 
-- LongRes(771) <= sub_result;
        -- when "0011111010" => 
-- LongRes(770) <= sub_result;
        -- when "0011111011" => 
-- LongRes(769) <= sub_result;
        -- when "0011111100" => 
-- LongRes(768) <= sub_result;
        -- when "0011111101" => 
-- LongRes(767) <= sub_result;
        -- when "0011111110" => 
-- LongRes(766) <= sub_result;
        -- when "0011111111" => 
-- LongRes(765) <= sub_result;
        -- when "0100000000" => 
-- LongRes(764) <= sub_result;
        -- when "0100000001" => 
-- LongRes(763) <= sub_result;
        -- when "0100000010" => 
-- LongRes(762) <= sub_result;
        -- when "0100000011" => 
-- LongRes(761) <= sub_result;
        -- when "0100000100" => 
-- LongRes(760) <= sub_result;
        -- when "0100000101" => 
-- LongRes(759) <= sub_result;
        -- when "0100000110" => 
-- LongRes(758) <= sub_result;
        -- when "0100000111" => 
-- LongRes(757) <= sub_result;
        -- when "0100001000" => 
-- LongRes(756) <= sub_result;
        -- when "0100001001" => 
-- LongRes(755) <= sub_result;
        -- when "0100001010" => 
-- LongRes(754) <= sub_result;
        -- when "0100001011" => 
-- LongRes(753) <= sub_result;
        -- when "0100001100" => 
-- LongRes(752) <= sub_result;
        -- when "0100001101" => 
-- LongRes(751) <= sub_result;
        -- when "0100001110" => 
-- LongRes(750) <= sub_result;
        -- when "0100001111" => 
-- LongRes(749) <= sub_result;
        -- when "0100010000" => 
-- LongRes(748) <= sub_result;
        -- when "0100010001" => 
-- LongRes(747) <= sub_result;
        -- when "0100010010" => 
-- LongRes(746) <= sub_result;
        -- when "0100010011" => 
-- LongRes(745) <= sub_result;
        -- when "0100010100" => 
-- LongRes(744) <= sub_result;
        -- when "0100010101" => 
-- LongRes(743) <= sub_result;
        -- when "0100010110" => 
-- LongRes(742) <= sub_result;
        -- when "0100010111" => 
-- LongRes(741) <= sub_result;
        -- when "0100011000" => 
-- LongRes(740) <= sub_result;
        -- when "0100011001" => 
-- LongRes(739) <= sub_result;
        -- when "0100011010" => 
-- LongRes(738) <= sub_result;
        -- when "0100011011" => 
-- LongRes(737) <= sub_result;
        -- when "0100011100" => 
-- LongRes(736) <= sub_result;
        -- when "0100011101" => 
-- LongRes(735) <= sub_result;
        -- when "0100011110" => 
-- LongRes(734) <= sub_result;
        -- when "0100011111" => 
-- LongRes(733) <= sub_result;
        -- when "0100100000" => 
-- LongRes(732) <= sub_result;
        -- when "0100100001" => 
-- LongRes(731) <= sub_result;
        -- when "0100100010" => 
-- LongRes(730) <= sub_result;
        -- when "0100100011" => 
-- LongRes(729) <= sub_result;
        -- when "0100100100" => 
-- LongRes(728) <= sub_result;
        -- when "0100100101" => 
-- LongRes(727) <= sub_result;
        -- when "0100100110" => 
-- LongRes(726) <= sub_result;
        -- when "0100100111" => 
-- LongRes(725) <= sub_result;
        -- when "0100101000" => 
-- LongRes(724) <= sub_result;
        -- when "0100101001" => 
-- LongRes(723) <= sub_result;
        -- when "0100101010" => 
-- LongRes(722) <= sub_result;
        -- when "0100101011" => 
-- LongRes(721) <= sub_result;
        -- when "0100101100" => 
-- LongRes(720) <= sub_result;
        -- when "0100101101" => 
-- LongRes(719) <= sub_result;
        -- when "0100101110" => 
-- LongRes(718) <= sub_result;
        -- when "0100101111" => 
-- LongRes(717) <= sub_result;
        -- when "0100110000" => 
-- LongRes(716) <= sub_result;
        -- when "0100110001" => 
-- LongRes(715) <= sub_result;
        -- when "0100110010" => 
-- LongRes(714) <= sub_result;
        -- when "0100110011" => 
-- LongRes(713) <= sub_result;
        -- when "0100110100" => 
-- LongRes(712) <= sub_result;
        -- when "0100110101" => 
-- LongRes(711) <= sub_result;
        -- when "0100110110" => 
-- LongRes(710) <= sub_result;
        -- when "0100110111" => 
-- LongRes(709) <= sub_result;
        -- when "0100111000" => 
-- LongRes(708) <= sub_result;
        -- when "0100111001" => 
-- LongRes(707) <= sub_result;
        -- when "0100111010" => 
-- LongRes(706) <= sub_result;
        -- when "0100111011" => 
-- LongRes(705) <= sub_result;
        -- when "0100111100" => 
-- LongRes(704) <= sub_result;
        -- when "0100111101" => 
-- LongRes(703) <= sub_result;
        -- when "0100111110" => 
-- LongRes(702) <= sub_result;
        -- when "0100111111" => 
-- LongRes(701) <= sub_result;
        -- when "0101000000" => 
-- LongRes(700) <= sub_result;
        -- when "0101000001" => 
-- LongRes(699) <= sub_result;
        -- when "0101000010" => 
-- LongRes(698) <= sub_result;
        -- when "0101000011" => 
-- LongRes(697) <= sub_result;
        -- when "0101000100" => 
-- LongRes(696) <= sub_result;
        -- when "0101000101" => 
-- LongRes(695) <= sub_result;
        -- when "0101000110" => 
-- LongRes(694) <= sub_result;
        -- when "0101000111" => 
-- LongRes(693) <= sub_result;
        -- when "0101001000" => 
-- LongRes(692) <= sub_result;
        -- when "0101001001" => 
-- LongRes(691) <= sub_result;
        -- when "0101001010" => 
-- LongRes(690) <= sub_result;
        -- when "0101001011" => 
-- LongRes(689) <= sub_result;
        -- when "0101001100" => 
-- LongRes(688) <= sub_result;
        -- when "0101001101" => 
-- LongRes(687) <= sub_result;
        -- when "0101001110" => 
-- LongRes(686) <= sub_result;
        -- when "0101001111" => 
-- LongRes(685) <= sub_result;
        -- when "0101010000" => 
-- LongRes(684) <= sub_result;
        -- when "0101010001" => 
-- LongRes(683) <= sub_result;
        -- when "0101010010" => 
-- LongRes(682) <= sub_result;
        -- when "0101010011" => 
-- LongRes(681) <= sub_result;
        -- when "0101010100" => 
-- LongRes(680) <= sub_result;
        -- when "0101010101" => 
-- LongRes(679) <= sub_result;
        -- when "0101010110" => 
-- LongRes(678) <= sub_result;
        -- when "0101010111" => 
-- LongRes(677) <= sub_result;
        -- when "0101011000" => 
-- LongRes(676) <= sub_result;
        -- when "0101011001" => 
-- LongRes(675) <= sub_result;
        -- when "0101011010" => 
-- LongRes(674) <= sub_result;
        -- when "0101011011" => 
-- LongRes(673) <= sub_result;
        -- when "0101011100" => 
-- LongRes(672) <= sub_result;
        -- when "0101011101" => 
-- LongRes(671) <= sub_result;
        -- when "0101011110" => 
-- LongRes(670) <= sub_result;
        -- when "0101011111" => 
-- LongRes(669) <= sub_result;
        -- when "0101100000" => 
-- LongRes(668) <= sub_result;
        -- when "0101100001" => 
-- LongRes(667) <= sub_result;
        -- when "0101100010" => 
-- LongRes(666) <= sub_result;
        -- when "0101100011" => 
-- LongRes(665) <= sub_result;
        -- when "0101100100" => 
-- LongRes(664) <= sub_result;
        -- when "0101100101" => 
-- LongRes(663) <= sub_result;
        -- when "0101100110" => 
-- LongRes(662) <= sub_result;
        -- when "0101100111" => 
-- LongRes(661) <= sub_result;
        -- when "0101101000" => 
-- LongRes(660) <= sub_result;
        -- when "0101101001" => 
-- LongRes(659) <= sub_result;
        -- when "0101101010" => 
-- LongRes(658) <= sub_result;
        -- when "0101101011" => 
-- LongRes(657) <= sub_result;
        -- when "0101101100" => 
-- LongRes(656) <= sub_result;
        -- when "0101101101" => 
-- LongRes(655) <= sub_result;
        -- when "0101101110" => 
-- LongRes(654) <= sub_result;
        -- when "0101101111" => 
-- LongRes(653) <= sub_result;
        -- when "0101110000" => 
-- LongRes(652) <= sub_result;
        -- when "0101110001" => 
-- LongRes(651) <= sub_result;
        -- when "0101110010" => 
-- LongRes(650) <= sub_result;
        -- when "0101110011" => 
-- LongRes(649) <= sub_result;
        -- when "0101110100" => 
-- LongRes(648) <= sub_result;
        -- when "0101110101" => 
-- LongRes(647) <= sub_result;
        -- when "0101110110" => 
-- LongRes(646) <= sub_result;
        -- when "0101110111" => 
-- LongRes(645) <= sub_result;
        -- when "0101111000" => 
-- LongRes(644) <= sub_result;
        -- when "0101111001" => 
-- LongRes(643) <= sub_result;
        -- when "0101111010" => 
-- LongRes(642) <= sub_result;
        -- when "0101111011" => 
-- LongRes(641) <= sub_result;
        -- when "0101111100" => 
-- LongRes(640) <= sub_result;
        -- when "0101111101" => 
-- LongRes(639) <= sub_result;
        -- when "0101111110" => 
-- LongRes(638) <= sub_result;
        -- when "0101111111" => 
-- LongRes(637) <= sub_result;
        -- when "0110000000" => 
-- LongRes(636) <= sub_result;
        -- when "0110000001" => 
-- LongRes(635) <= sub_result;
        -- when "0110000010" => 
-- LongRes(634) <= sub_result;
        -- when "0110000011" => 
-- LongRes(633) <= sub_result;
        -- when "0110000100" => 
-- LongRes(632) <= sub_result;
        -- when "0110000101" => 
-- LongRes(631) <= sub_result;
        -- when "0110000110" => 
-- LongRes(630) <= sub_result;
        -- when "0110000111" => 
-- LongRes(629) <= sub_result;
        -- when "0110001000" => 
-- LongRes(628) <= sub_result;
        -- when "0110001001" => 
-- LongRes(627) <= sub_result;
        -- when "0110001010" => 
-- LongRes(626) <= sub_result;
        -- when "0110001011" => 
-- LongRes(625) <= sub_result;
        -- when "0110001100" => 
-- LongRes(624) <= sub_result;
        -- when "0110001101" => 
-- LongRes(623) <= sub_result;
        -- when "0110001110" => 
-- LongRes(622) <= sub_result;
        -- when "0110001111" => 
-- LongRes(621) <= sub_result;
        -- when "0110010000" => 
-- LongRes(620) <= sub_result;
        -- when "0110010001" => 
-- LongRes(619) <= sub_result;
        -- when "0110010010" => 
-- LongRes(618) <= sub_result;
        -- when "0110010011" => 
-- LongRes(617) <= sub_result;
        -- when "0110010100" => 
-- LongRes(616) <= sub_result;
        -- when "0110010101" => 
-- LongRes(615) <= sub_result;
        -- when "0110010110" => 
-- LongRes(614) <= sub_result;
        -- when "0110010111" => 
-- LongRes(613) <= sub_result;
        -- when "0110011000" => 
-- LongRes(612) <= sub_result;
        -- when "0110011001" => 
-- LongRes(611) <= sub_result;
        -- when "0110011010" => 
-- LongRes(610) <= sub_result;
        -- when "0110011011" => 
-- LongRes(609) <= sub_result;
        -- when "0110011100" => 
-- LongRes(608) <= sub_result;
        -- when "0110011101" => 
-- LongRes(607) <= sub_result;
        -- when "0110011110" => 
-- LongRes(606) <= sub_result;
        -- when "0110011111" => 
-- LongRes(605) <= sub_result;
        -- when "0110100000" => 
-- LongRes(604) <= sub_result;
        -- when "0110100001" => 
-- LongRes(603) <= sub_result;
        -- when "0110100010" => 
-- LongRes(602) <= sub_result;
        -- when "0110100011" => 
-- LongRes(601) <= sub_result;
        -- when "0110100100" => 
-- LongRes(600) <= sub_result;
        -- when "0110100101" => 
-- LongRes(599) <= sub_result;
        -- when "0110100110" => 
-- LongRes(598) <= sub_result;
        -- when "0110100111" => 
-- LongRes(597) <= sub_result;
        -- when "0110101000" => 
-- LongRes(596) <= sub_result;
        -- when "0110101001" => 
-- LongRes(595) <= sub_result;
        -- when "0110101010" => 
-- LongRes(594) <= sub_result;
        -- when "0110101011" => 
-- LongRes(593) <= sub_result;
        -- when "0110101100" => 
-- LongRes(592) <= sub_result;
        -- when "0110101101" => 
-- LongRes(591) <= sub_result;
        -- when "0110101110" => 
-- LongRes(590) <= sub_result;
        -- when "0110101111" => 
-- LongRes(589) <= sub_result;
        -- when "0110110000" => 
-- LongRes(588) <= sub_result;
        -- when "0110110001" => 
-- LongRes(587) <= sub_result;
        -- when "0110110010" => 
-- LongRes(586) <= sub_result;
        -- when "0110110011" => 
-- LongRes(585) <= sub_result;
        -- when "0110110100" => 
-- LongRes(584) <= sub_result;
        -- when "0110110101" => 
-- LongRes(583) <= sub_result;
        -- when "0110110110" => 
-- LongRes(582) <= sub_result;
        -- when "0110110111" => 
-- LongRes(581) <= sub_result;
        -- when "0110111000" => 
-- LongRes(580) <= sub_result;
        -- when "0110111001" => 
-- LongRes(579) <= sub_result;
        -- when "0110111010" => 
-- LongRes(578) <= sub_result;
        -- when "0110111011" => 
-- LongRes(577) <= sub_result;
        -- when "0110111100" => 
-- LongRes(576) <= sub_result;
        -- when "0110111101" => 
-- LongRes(575) <= sub_result;
        -- when "0110111110" => 
-- LongRes(574) <= sub_result;
        -- when "0110111111" => 
-- LongRes(573) <= sub_result;
        -- when "0111000000" => 
-- LongRes(572) <= sub_result;
        -- when "0111000001" => 
-- LongRes(571) <= sub_result;
        -- when "0111000010" => 
-- LongRes(570) <= sub_result;
        -- when "0111000011" => 
-- LongRes(569) <= sub_result;
        -- when "0111000100" => 
-- LongRes(568) <= sub_result;
        -- when "0111000101" => 
-- LongRes(567) <= sub_result;
        -- when "0111000110" => 
-- LongRes(566) <= sub_result;
        -- when "0111000111" => 
-- LongRes(565) <= sub_result;
        -- when "0111001000" => 
-- LongRes(564) <= sub_result;
        -- when "0111001001" => 
-- LongRes(563) <= sub_result;
        -- when "0111001010" => 
-- LongRes(562) <= sub_result;
        -- when "0111001011" => 
-- LongRes(561) <= sub_result;
        -- when "0111001100" => 
-- LongRes(560) <= sub_result;
        -- when "0111001101" => 
-- LongRes(559) <= sub_result;
        -- when "0111001110" => 
-- LongRes(558) <= sub_result;
        -- when "0111001111" => 
-- LongRes(557) <= sub_result;
        -- when "0111010000" => 
-- LongRes(556) <= sub_result;
        -- when "0111010001" => 
-- LongRes(555) <= sub_result;
        -- when "0111010010" => 
-- LongRes(554) <= sub_result;
        -- when "0111010011" => 
-- LongRes(553) <= sub_result;
        -- when "0111010100" => 
-- LongRes(552) <= sub_result;
        -- when "0111010101" => 
-- LongRes(551) <= sub_result;
        -- when "0111010110" => 
-- LongRes(550) <= sub_result;
        -- when "0111010111" => 
-- LongRes(549) <= sub_result;
        -- when "0111011000" => 
-- LongRes(548) <= sub_result;
        -- when "0111011001" => 
-- LongRes(547) <= sub_result;
        -- when "0111011010" => 
-- LongRes(546) <= sub_result;
        -- when "0111011011" => 
-- LongRes(545) <= sub_result;
        -- when "0111011100" => 
-- LongRes(544) <= sub_result;
        -- when "0111011101" => 
-- LongRes(543) <= sub_result;
        -- when "0111011110" => 
-- LongRes(542) <= sub_result;
        -- when "0111011111" => 
-- LongRes(541) <= sub_result;
        -- when "0111100000" => 
-- LongRes(540) <= sub_result;
        -- when "0111100001" => 
-- LongRes(539) <= sub_result;
        -- when "0111100010" => 
-- LongRes(538) <= sub_result;
        -- when "0111100011" => 
-- LongRes(537) <= sub_result;
        -- when "0111100100" => 
-- LongRes(536) <= sub_result;
        -- when "0111100101" => 
-- LongRes(535) <= sub_result;
        -- when "0111100110" => 
-- LongRes(534) <= sub_result;
        -- when "0111100111" => 
-- LongRes(533) <= sub_result;
        -- when "0111101000" => 
-- LongRes(532) <= sub_result;
        -- when "0111101001" => 
-- LongRes(531) <= sub_result;
        -- when "0111101010" => 
-- LongRes(530) <= sub_result;
        -- when "0111101011" => 
-- LongRes(529) <= sub_result;
        -- when "0111101100" => 
-- LongRes(528) <= sub_result;
        -- when "0111101101" => 
-- LongRes(527) <= sub_result;
        -- when "0111101110" => 
-- LongRes(526) <= sub_result;
        -- when "0111101111" => 
-- LongRes(525) <= sub_result;
        -- when "0111110000" => 
-- LongRes(524) <= sub_result;
        -- when "0111110001" => 
-- LongRes(523) <= sub_result;
        -- when "0111110010" => 
-- LongRes(522) <= sub_result;
        -- when "0111110011" => 
-- LongRes(521) <= sub_result;
        -- when "0111110100" => 
-- LongRes(520) <= sub_result;
        -- when "0111110101" => 
-- LongRes(519) <= sub_result;
        -- when "0111110110" => 
-- LongRes(518) <= sub_result;
        -- when "0111110111" => 
-- LongRes(517) <= sub_result;
        -- when "0111111000" => 
-- LongRes(516) <= sub_result;
        -- when "0111111001" => 
-- LongRes(515) <= sub_result;
        -- when "0111111010" => 
-- LongRes(514) <= sub_result;
        -- when "0111111011" => 
-- LongRes(513) <= sub_result;
        -- when "0111111100" => 
-- LongRes(512) <= sub_result;
        -- when "0111111101" => 
-- LongRes(511) <= sub_result;
        -- when "0111111110" => 
-- LongRes(510) <= sub_result;
        -- when "0111111111" => 
-- LongRes(509) <= sub_result;
        -- when "1000000000" => 
-- LongRes(508) <= sub_result;
        -- when "1000000001" => 
-- LongRes(507) <= sub_result;
        -- when "1000000010" => 
-- LongRes(506) <= sub_result;
        -- when "1000000011" => 
-- LongRes(505) <= sub_result;
        -- when "1000000100" => 
-- LongRes(504) <= sub_result;
        -- when "1000000101" => 
-- LongRes(503) <= sub_result;
        -- when "1000000110" => 
-- LongRes(502) <= sub_result;
        -- when "1000000111" => 
-- LongRes(501) <= sub_result;
        -- when "1000001000" => 
-- LongRes(500) <= sub_result;
        -- when "1000001001" => 
-- LongRes(499) <= sub_result;
        -- when "1000001010" => 
-- LongRes(498) <= sub_result;
        -- when "1000001011" => 
-- LongRes(497) <= sub_result;
        -- when "1000001100" => 
-- LongRes(496) <= sub_result;
        -- when "1000001101" => 
-- LongRes(495) <= sub_result;
        -- when "1000001110" => 
-- LongRes(494) <= sub_result;
        -- when "1000001111" => 
-- LongRes(493) <= sub_result;
        -- when "1000010000" => 
-- LongRes(492) <= sub_result;
        -- when "1000010001" => 
-- LongRes(491) <= sub_result;
        -- when "1000010010" => 
-- LongRes(490) <= sub_result;
        -- when "1000010011" => 
-- LongRes(489) <= sub_result;
        -- when "1000010100" => 
-- LongRes(488) <= sub_result;
        -- when "1000010101" => 
-- LongRes(487) <= sub_result;
        -- when "1000010110" => 
-- LongRes(486) <= sub_result;
        -- when "1000010111" => 
-- LongRes(485) <= sub_result;
        -- when "1000011000" => 
-- LongRes(484) <= sub_result;
        -- when "1000011001" => 
-- LongRes(483) <= sub_result;
        -- when "1000011010" => 
-- LongRes(482) <= sub_result;
        -- when "1000011011" => 
-- LongRes(481) <= sub_result;
        -- when "1000011100" => 
-- LongRes(480) <= sub_result;
        -- when "1000011101" => 
-- LongRes(479) <= sub_result;
        -- when "1000011110" => 
-- LongRes(478) <= sub_result;
        -- when "1000011111" => 
-- LongRes(477) <= sub_result;
        -- when "1000100000" => 
-- LongRes(476) <= sub_result;
        -- when "1000100001" => 
-- LongRes(475) <= sub_result;
        -- when "1000100010" => 
-- LongRes(474) <= sub_result;
        -- when "1000100011" => 
-- LongRes(473) <= sub_result;
        -- when "1000100100" => 
-- LongRes(472) <= sub_result;
        -- when "1000100101" => 
-- LongRes(471) <= sub_result;
        -- when "1000100110" => 
-- LongRes(470) <= sub_result;
        -- when "1000100111" => 
-- LongRes(469) <= sub_result;
        -- when "1000101000" => 
-- LongRes(468) <= sub_result;
        -- when "1000101001" => 
-- LongRes(467) <= sub_result;
        -- when "1000101010" => 
-- LongRes(466) <= sub_result;
        -- when "1000101011" => 
-- LongRes(465) <= sub_result;
        -- when "1000101100" => 
-- LongRes(464) <= sub_result;
        -- when "1000101101" => 
-- LongRes(463) <= sub_result;
        -- when "1000101110" => 
-- LongRes(462) <= sub_result;
        -- when "1000101111" => 
-- LongRes(461) <= sub_result;
        -- when "1000110000" => 
-- LongRes(460) <= sub_result;
        -- when "1000110001" => 
-- LongRes(459) <= sub_result;
        -- when "1000110010" => 
-- LongRes(458) <= sub_result;
        -- when "1000110011" => 
-- LongRes(457) <= sub_result;
        -- when "1000110100" => 
-- LongRes(456) <= sub_result;
        -- when "1000110101" => 
-- LongRes(455) <= sub_result;
        -- when "1000110110" => 
-- LongRes(454) <= sub_result;
        -- when "1000110111" => 
-- LongRes(453) <= sub_result;
        -- when "1000111000" => 
-- LongRes(452) <= sub_result;
        -- when "1000111001" => 
-- LongRes(451) <= sub_result;
        -- when "1000111010" => 
-- LongRes(450) <= sub_result;
        -- when "1000111011" => 
-- LongRes(449) <= sub_result;
        -- when "1000111100" => 
-- LongRes(448) <= sub_result;
        -- when "1000111101" => 
-- LongRes(447) <= sub_result;
        -- when "1000111110" => 
-- LongRes(446) <= sub_result;
        -- when "1000111111" => 
-- LongRes(445) <= sub_result;
        -- when "1001000000" => 
-- LongRes(444) <= sub_result;
        -- when "1001000001" => 
-- LongRes(443) <= sub_result;
        -- when "1001000010" => 
-- LongRes(442) <= sub_result;
        -- when "1001000011" => 
-- LongRes(441) <= sub_result;
        -- when "1001000100" => 
-- LongRes(440) <= sub_result;
        -- when "1001000101" => 
-- LongRes(439) <= sub_result;
        -- when "1001000110" => 
-- LongRes(438) <= sub_result;
        -- when "1001000111" => 
-- LongRes(437) <= sub_result;
        -- when "1001001000" => 
-- LongRes(436) <= sub_result;
        -- when "1001001001" => 
-- LongRes(435) <= sub_result;
        -- when "1001001010" => 
-- LongRes(434) <= sub_result;
        -- when "1001001011" => 
-- LongRes(433) <= sub_result;
        -- when "1001001100" => 
-- LongRes(432) <= sub_result;
        -- when "1001001101" => 
-- LongRes(431) <= sub_result;
        -- when "1001001110" => 
-- LongRes(430) <= sub_result;
        -- when "1001001111" => 
-- LongRes(429) <= sub_result;
        -- when "1001010000" => 
-- LongRes(428) <= sub_result;
        -- when "1001010001" => 
-- LongRes(427) <= sub_result;
        -- when "1001010010" => 
-- LongRes(426) <= sub_result;
        -- when "1001010011" => 
-- LongRes(425) <= sub_result;
        -- when "1001010100" => 
-- LongRes(424) <= sub_result;
        -- when "1001010101" => 
-- LongRes(423) <= sub_result;
        -- when "1001010110" => 
-- LongRes(422) <= sub_result;
        -- when "1001010111" => 
-- LongRes(421) <= sub_result;
        -- when "1001011000" => 
-- LongRes(420) <= sub_result;
        -- when "1001011001" => 
-- LongRes(419) <= sub_result;
        -- when "1001011010" => 
-- LongRes(418) <= sub_result;
        -- when "1001011011" => 
-- LongRes(417) <= sub_result;
        -- when "1001011100" => 
-- LongRes(416) <= sub_result;
        -- when "1001011101" => 
-- LongRes(415) <= sub_result;
        -- when "1001011110" => 
-- LongRes(414) <= sub_result;
        -- when "1001011111" => 
-- LongRes(413) <= sub_result;
        -- when "1001100000" => 
-- LongRes(412) <= sub_result;
        -- when "1001100001" => 
-- LongRes(411) <= sub_result;
        -- when "1001100010" => 
-- LongRes(410) <= sub_result;
        -- when "1001100011" => 
-- LongRes(409) <= sub_result;
        -- when "1001100100" => 
-- LongRes(408) <= sub_result;
        -- when "1001100101" => 
-- LongRes(407) <= sub_result;
        -- when "1001100110" => 
-- LongRes(406) <= sub_result;
        -- when "1001100111" => 
-- LongRes(405) <= sub_result;
        -- when "1001101000" => 
-- LongRes(404) <= sub_result;
        -- when "1001101001" => 
-- LongRes(403) <= sub_result;
        -- when "1001101010" => 
-- LongRes(402) <= sub_result;
        -- when "1001101011" => 
-- LongRes(401) <= sub_result;
        -- when "1001101100" => 
-- LongRes(400) <= sub_result;
        -- when "1001101101" => 
-- LongRes(399) <= sub_result;
        -- when "1001101110" => 
-- LongRes(398) <= sub_result;
        -- when "1001101111" => 
-- LongRes(397) <= sub_result;
        -- when "1001110000" => 
-- LongRes(396) <= sub_result;
        -- when "1001110001" => 
-- LongRes(395) <= sub_result;
        -- when "1001110010" => 
-- LongRes(394) <= sub_result;
        -- when "1001110011" => 
-- LongRes(393) <= sub_result;
        -- when "1001110100" => 
-- LongRes(392) <= sub_result;
        -- when "1001110101" => 
-- LongRes(391) <= sub_result;
        -- when "1001110110" => 
-- LongRes(390) <= sub_result;
        -- when "1001110111" => 
-- LongRes(389) <= sub_result;
        -- when "1001111000" => 
-- LongRes(388) <= sub_result;
        -- when "1001111001" => 
-- LongRes(387) <= sub_result;
        -- when "1001111010" => 
-- LongRes(386) <= sub_result;
        -- when "1001111011" => 
-- LongRes(385) <= sub_result;
        -- when "1001111100" => 
-- LongRes(384) <= sub_result;
        -- when "1001111101" => 
-- LongRes(383) <= sub_result;
        -- when "1001111110" => 
-- LongRes(382) <= sub_result;
        -- when "1001111111" => 
-- LongRes(381) <= sub_result;
        -- when "1010000000" => 
-- LongRes(380) <= sub_result;
        -- when "1010000001" => 
-- LongRes(379) <= sub_result;
        -- when "1010000010" => 
-- LongRes(378) <= sub_result;
        -- when "1010000011" => 
-- LongRes(377) <= sub_result;
        -- when "1010000100" => 
-- LongRes(376) <= sub_result;
        -- when "1010000101" => 
-- LongRes(375) <= sub_result;
        -- when "1010000110" => 
-- LongRes(374) <= sub_result;
        -- when "1010000111" => 
-- LongRes(373) <= sub_result;
        -- when "1010001000" => 
-- LongRes(372) <= sub_result;
        -- when "1010001001" => 
-- LongRes(371) <= sub_result;
        -- when "1010001010" => 
-- LongRes(370) <= sub_result;
        -- when "1010001011" => 
-- LongRes(369) <= sub_result;
        -- when "1010001100" => 
-- LongRes(368) <= sub_result;
        -- when "1010001101" => 
-- LongRes(367) <= sub_result;
        -- when "1010001110" => 
-- LongRes(366) <= sub_result;
        -- when "1010001111" => 
-- LongRes(365) <= sub_result;
        -- when "1010010000" => 
-- LongRes(364) <= sub_result;
        -- when "1010010001" => 
-- LongRes(363) <= sub_result;
        -- when "1010010010" => 
-- LongRes(362) <= sub_result;
        -- when "1010010011" => 
-- LongRes(361) <= sub_result;
        -- when "1010010100" => 
-- LongRes(360) <= sub_result;
        -- when "1010010101" => 
-- LongRes(359) <= sub_result;
        -- when "1010010110" => 
-- LongRes(358) <= sub_result;
        -- when "1010010111" => 
-- LongRes(357) <= sub_result;
        -- when "1010011000" => 
-- LongRes(356) <= sub_result;
        -- when "1010011001" => 
-- LongRes(355) <= sub_result;
        -- when "1010011010" => 
-- LongRes(354) <= sub_result;
        -- when "1010011011" => 
-- LongRes(353) <= sub_result;
        -- when "1010011100" => 
-- LongRes(352) <= sub_result;
        -- when "1010011101" => 
-- LongRes(351) <= sub_result;
        -- when "1010011110" => 
-- LongRes(350) <= sub_result;
        -- when "1010011111" => 
-- LongRes(349) <= sub_result;
        -- when "1010100000" => 
-- LongRes(348) <= sub_result;
        -- when "1010100001" => 
-- LongRes(347) <= sub_result;
        -- when "1010100010" => 
-- LongRes(346) <= sub_result;
        -- when "1010100011" => 
-- LongRes(345) <= sub_result;
        -- when "1010100100" => 
-- LongRes(344) <= sub_result;
        -- when "1010100101" => 
-- LongRes(343) <= sub_result;
        -- when "1010100110" => 
-- LongRes(342) <= sub_result;
        -- when "1010100111" => 
-- LongRes(341) <= sub_result;
        -- when "1010101000" => 
-- LongRes(340) <= sub_result;
        -- when "1010101001" => 
-- LongRes(339) <= sub_result;
        -- when "1010101010" => 
-- LongRes(338) <= sub_result;
        -- when "1010101011" => 
-- LongRes(337) <= sub_result;
        -- when "1010101100" => 
-- LongRes(336) <= sub_result;
        -- when "1010101101" => 
-- LongRes(335) <= sub_result;
        -- when "1010101110" => 
-- LongRes(334) <= sub_result;
        -- when "1010101111" => 
-- LongRes(333) <= sub_result;
        -- when "1010110000" => 
-- LongRes(332) <= sub_result;
        -- when "1010110001" => 
-- LongRes(331) <= sub_result;
        -- when "1010110010" => 
-- LongRes(330) <= sub_result;
        -- when "1010110011" => 
-- LongRes(329) <= sub_result;
        -- when "1010110100" => 
-- LongRes(328) <= sub_result;
        -- when "1010110101" => 
-- LongRes(327) <= sub_result;
        -- when "1010110110" => 
-- LongRes(326) <= sub_result;
        -- when "1010110111" => 
-- LongRes(325) <= sub_result;
        -- when "1010111000" => 
-- LongRes(324) <= sub_result;
        -- when "1010111001" => 
-- LongRes(323) <= sub_result;
        -- when "1010111010" => 
-- LongRes(322) <= sub_result;
        -- when "1010111011" => 
-- LongRes(321) <= sub_result;
        -- when "1010111100" => 
-- LongRes(320) <= sub_result;
        -- when "1010111101" => 
-- LongRes(319) <= sub_result;
        -- when "1010111110" => 
-- LongRes(318) <= sub_result;
        -- when "1010111111" => 
-- LongRes(317) <= sub_result;
        -- when "1011000000" => 
-- LongRes(316) <= sub_result;
        -- when "1011000001" => 
-- LongRes(315) <= sub_result;
        -- when "1011000010" => 
-- LongRes(314) <= sub_result;
        -- when "1011000011" => 
-- LongRes(313) <= sub_result;
        -- when "1011000100" => 
-- LongRes(312) <= sub_result;
        -- when "1011000101" => 
-- LongRes(311) <= sub_result;
        -- when "1011000110" => 
-- LongRes(310) <= sub_result;
        -- when "1011000111" => 
-- LongRes(309) <= sub_result;
        -- when "1011001000" => 
-- LongRes(308) <= sub_result;
        -- when "1011001001" => 
-- LongRes(307) <= sub_result;
        -- when "1011001010" => 
-- LongRes(306) <= sub_result;
        -- when "1011001011" => 
-- LongRes(305) <= sub_result;
        -- when "1011001100" => 
-- LongRes(304) <= sub_result;
        -- when "1011001101" => 
-- LongRes(303) <= sub_result;
        -- when "1011001110" => 
-- LongRes(302) <= sub_result;
        -- when "1011001111" => 
-- LongRes(301) <= sub_result;
        -- when "1011010000" => 
-- LongRes(300) <= sub_result;
        -- when "1011010001" => 
-- LongRes(299) <= sub_result;
        -- when "1011010010" => 
-- LongRes(298) <= sub_result;
        -- when "1011010011" => 
-- LongRes(297) <= sub_result;
        -- when "1011010100" => 
-- LongRes(296) <= sub_result;
        -- when "1011010101" => 
-- LongRes(295) <= sub_result;
        -- when "1011010110" => 
-- LongRes(294) <= sub_result;
        -- when "1011010111" => 
-- LongRes(293) <= sub_result;
        -- when "1011011000" => 
-- LongRes(292) <= sub_result;
        -- when "1011011001" => 
-- LongRes(291) <= sub_result;
        -- when "1011011010" => 
-- LongRes(290) <= sub_result;
        -- when "1011011011" => 
-- LongRes(289) <= sub_result;
        -- when "1011011100" => 
-- LongRes(288) <= sub_result;
        -- when "1011011101" => 
-- LongRes(287) <= sub_result;
        -- when "1011011110" => 
-- LongRes(286) <= sub_result;
        -- when "1011011111" => 
-- LongRes(285) <= sub_result;
        -- when "1011100000" => 
-- LongRes(284) <= sub_result;
        -- when "1011100001" => 
-- LongRes(283) <= sub_result;
        -- when "1011100010" => 
-- LongRes(282) <= sub_result;
        -- when "1011100011" => 
-- LongRes(281) <= sub_result;
        -- when "1011100100" => 
-- LongRes(280) <= sub_result;
        -- when "1011100101" => 
-- LongRes(279) <= sub_result;
        -- when "1011100110" => 
-- LongRes(278) <= sub_result;
        -- when "1011100111" => 
-- LongRes(277) <= sub_result;
        -- when "1011101000" => 
-- LongRes(276) <= sub_result;
        -- when "1011101001" => 
-- LongRes(275) <= sub_result;
        -- when "1011101010" => 
-- LongRes(274) <= sub_result;
        -- when "1011101011" => 
-- LongRes(273) <= sub_result;
        -- when "1011101100" => 
-- LongRes(272) <= sub_result;
        -- when "1011101101" => 
-- LongRes(271) <= sub_result;
        -- when "1011101110" => 
-- LongRes(270) <= sub_result;
        -- when "1011101111" => 
-- LongRes(269) <= sub_result;
        -- when "1011110000" => 
-- LongRes(268) <= sub_result;
        -- when "1011110001" => 
-- LongRes(267) <= sub_result;
        -- when "1011110010" => 
-- LongRes(266) <= sub_result;
        -- when "1011110011" => 
-- LongRes(265) <= sub_result;
        -- when "1011110100" => 
-- LongRes(264) <= sub_result;
        -- when "1011110101" => 
-- LongRes(263) <= sub_result;
        -- when "1011110110" => 
-- LongRes(262) <= sub_result;
        -- when "1011110111" => 
-- LongRes(261) <= sub_result;
        -- when "1011111000" => 
-- LongRes(260) <= sub_result;
        -- when "1011111001" => 
-- LongRes(259) <= sub_result;
        -- when "1011111010" => 
-- LongRes(258) <= sub_result;
        -- when "1011111011" => 
-- LongRes(257) <= sub_result;
        -- when "1011111100" => 
-- LongRes(256) <= sub_result;
        -- when "1011111101" => 
-- LongRes(255) <= sub_result;
        -- when "1011111110" => 
-- LongRes(254) <= sub_result;
        -- when "1011111111" => 
-- LongRes(253) <= sub_result;
        -- when "1100000000" => 
-- LongRes(252) <= sub_result;
        -- when "1100000001" => 
-- LongRes(251) <= sub_result;
        -- when "1100000010" => 
-- LongRes(250) <= sub_result;
        -- when "1100000011" => 
-- LongRes(249) <= sub_result;
        -- when "1100000100" => 
-- LongRes(248) <= sub_result;
        -- when "1100000101" => 
-- LongRes(247) <= sub_result;
        -- when "1100000110" => 
-- LongRes(246) <= sub_result;
        -- when "1100000111" => 
-- LongRes(245) <= sub_result;
        -- when "1100001000" => 
-- LongRes(244) <= sub_result;
        -- when "1100001001" => 
-- LongRes(243) <= sub_result;
        -- when "1100001010" => 
-- LongRes(242) <= sub_result;
        -- when "1100001011" => 
-- LongRes(241) <= sub_result;
        -- when "1100001100" => 
-- LongRes(240) <= sub_result;
        -- when "1100001101" => 
-- LongRes(239) <= sub_result;
        -- when "1100001110" => 
-- LongRes(238) <= sub_result;
        -- when "1100001111" => 
-- LongRes(237) <= sub_result;
        -- when "1100010000" => 
-- LongRes(236) <= sub_result;
        -- when "1100010001" => 
-- LongRes(235) <= sub_result;
        -- when "1100010010" => 
-- LongRes(234) <= sub_result;
        -- when "1100010011" => 
-- LongRes(233) <= sub_result;
        -- when "1100010100" => 
-- LongRes(232) <= sub_result;
        -- when "1100010101" => 
-- LongRes(231) <= sub_result;
        -- when "1100010110" => 
-- LongRes(230) <= sub_result;
        -- when "1100010111" => 
-- LongRes(229) <= sub_result;
        -- when "1100011000" => 
-- LongRes(228) <= sub_result;
        -- when "1100011001" => 
-- LongRes(227) <= sub_result;
        -- when "1100011010" => 
-- LongRes(226) <= sub_result;
        -- when "1100011011" => 
-- LongRes(225) <= sub_result;
        -- when "1100011100" => 
-- LongRes(224) <= sub_result;
        -- when "1100011101" => 
-- LongRes(223) <= sub_result;
        -- when "1100011110" => 
-- LongRes(222) <= sub_result;
        -- when "1100011111" => 
-- LongRes(221) <= sub_result;
        -- when "1100100000" => 
-- LongRes(220) <= sub_result;
        -- when "1100100001" => 
-- LongRes(219) <= sub_result;
        -- when "1100100010" => 
-- LongRes(218) <= sub_result;
        -- when "1100100011" => 
-- LongRes(217) <= sub_result;
        -- when "1100100100" => 
-- LongRes(216) <= sub_result;
        -- when "1100100101" => 
-- LongRes(215) <= sub_result;
        -- when "1100100110" => 
-- LongRes(214) <= sub_result;
        -- when "1100100111" => 
-- LongRes(213) <= sub_result;
        -- when "1100101000" => 
-- LongRes(212) <= sub_result;
        -- when "1100101001" => 
-- LongRes(211) <= sub_result;
        -- when "1100101010" => 
-- LongRes(210) <= sub_result;
        -- when "1100101011" => 
-- LongRes(209) <= sub_result;
        -- when "1100101100" => 
-- LongRes(208) <= sub_result;
        -- when "1100101101" => 
-- LongRes(207) <= sub_result;
        -- when "1100101110" => 
-- LongRes(206) <= sub_result;
        -- when "1100101111" => 
-- LongRes(205) <= sub_result;
        -- when "1100110000" => 
-- LongRes(204) <= sub_result;
        -- when "1100110001" => 
-- LongRes(203) <= sub_result;
        -- when "1100110010" => 
-- LongRes(202) <= sub_result;
        -- when "1100110011" => 
-- LongRes(201) <= sub_result;
        -- when "1100110100" => 
-- LongRes(200) <= sub_result;
        -- when "1100110101" => 
-- LongRes(199) <= sub_result;
        -- when "1100110110" => 
-- LongRes(198) <= sub_result;
        -- when "1100110111" => 
-- LongRes(197) <= sub_result;
        -- when "1100111000" => 
-- LongRes(196) <= sub_result;
        -- when "1100111001" => 
-- LongRes(195) <= sub_result;
        -- when "1100111010" => 
-- LongRes(194) <= sub_result;
        -- when "1100111011" => 
-- LongRes(193) <= sub_result;
        -- when "1100111100" => 
-- LongRes(192) <= sub_result;
        -- when "1100111101" => 
-- LongRes(191) <= sub_result;
        -- when "1100111110" => 
-- LongRes(190) <= sub_result;
        -- when "1100111111" => 
-- LongRes(189) <= sub_result;
        -- when "1101000000" => 
-- LongRes(188) <= sub_result;
        -- when "1101000001" => 
-- LongRes(187) <= sub_result;
        -- when "1101000010" => 
-- LongRes(186) <= sub_result;
        -- when "1101000011" => 
-- LongRes(185) <= sub_result;
        -- when "1101000100" => 
-- LongRes(184) <= sub_result;
        -- when "1101000101" => 
-- LongRes(183) <= sub_result;
        -- when "1101000110" => 
-- LongRes(182) <= sub_result;
        -- when "1101000111" => 
-- LongRes(181) <= sub_result;
        -- when "1101001000" => 
-- LongRes(180) <= sub_result;
        -- when "1101001001" => 
-- LongRes(179) <= sub_result;
        -- when "1101001010" => 
-- LongRes(178) <= sub_result;
        -- when "1101001011" => 
-- LongRes(177) <= sub_result;
        -- when "1101001100" => 
-- LongRes(176) <= sub_result;
        -- when "1101001101" => 
-- LongRes(175) <= sub_result;
        -- when "1101001110" => 
-- LongRes(174) <= sub_result;
        -- when "1101001111" => 
-- LongRes(173) <= sub_result;
        -- when "1101010000" => 
-- LongRes(172) <= sub_result;
        -- when "1101010001" => 
-- LongRes(171) <= sub_result;
        -- when "1101010010" => 
-- LongRes(170) <= sub_result;
        -- when "1101010011" => 
-- LongRes(169) <= sub_result;
        -- when "1101010100" => 
-- LongRes(168) <= sub_result;
        -- when "1101010101" => 
-- LongRes(167) <= sub_result;
        -- when "1101010110" => 
-- LongRes(166) <= sub_result;
        -- when "1101010111" => 
-- LongRes(165) <= sub_result;
        -- when "1101011000" => 
-- LongRes(164) <= sub_result;
        -- when "1101011001" => 
-- LongRes(163) <= sub_result;
        -- when "1101011010" => 
-- LongRes(162) <= sub_result;
        -- when "1101011011" => 
-- LongRes(161) <= sub_result;
        -- when "1101011100" => 
-- LongRes(160) <= sub_result;
        -- when "1101011101" => 
-- LongRes(159) <= sub_result;
        -- when "1101011110" => 
-- LongRes(158) <= sub_result;
        -- when "1101011111" => 
-- LongRes(157) <= sub_result;
        -- when "1101100000" => 
-- LongRes(156) <= sub_result;
        -- when "1101100001" => 
-- LongRes(155) <= sub_result;
        -- when "1101100010" => 
-- LongRes(154) <= sub_result;
        -- when "1101100011" => 
-- LongRes(153) <= sub_result;
        -- when "1101100100" => 
-- LongRes(152) <= sub_result;
        -- when "1101100101" => 
-- LongRes(151) <= sub_result;
        -- when "1101100110" => 
-- LongRes(150) <= sub_result;
        -- when "1101100111" => 
-- LongRes(149) <= sub_result;
        -- when "1101101000" => 
-- LongRes(148) <= sub_result;
        -- when "1101101001" => 
-- LongRes(147) <= sub_result;
        -- when "1101101010" => 
-- LongRes(146) <= sub_result;
        -- when "1101101011" => 
-- LongRes(145) <= sub_result;
        -- when "1101101100" => 
-- LongRes(144) <= sub_result;
        -- when "1101101101" => 
-- LongRes(143) <= sub_result;
        -- when "1101101110" => 
-- LongRes(142) <= sub_result;
        -- when "1101101111" => 
-- LongRes(141) <= sub_result;
        -- when "1101110000" => 
-- LongRes(140) <= sub_result;
        -- when "1101110001" => 
-- LongRes(139) <= sub_result;
        -- when "1101110010" => 
-- LongRes(138) <= sub_result;
        -- when "1101110011" => 
-- LongRes(137) <= sub_result;
        -- when "1101110100" => 
-- LongRes(136) <= sub_result;
        -- when "1101110101" => 
-- LongRes(135) <= sub_result;
        -- when "1101110110" => 
-- LongRes(134) <= sub_result;
        -- when "1101110111" => 
-- LongRes(133) <= sub_result;
        -- when "1101111000" => 
-- LongRes(132) <= sub_result;
        -- when "1101111001" => 
-- LongRes(131) <= sub_result;
        -- when "1101111010" => 
-- LongRes(130) <= sub_result;
        -- when "1101111011" => 
-- LongRes(129) <= sub_result;
        -- when "1101111100" => 
-- LongRes(128) <= sub_result;
        -- when "1101111101" => 
-- LongRes(127) <= sub_result;
        -- when "1101111110" => 
-- LongRes(126) <= sub_result;
        -- when "1101111111" => 
-- LongRes(125) <= sub_result;
        -- when "1110000000" => 
-- LongRes(124) <= sub_result;
        -- when "1110000001" => 
-- LongRes(123) <= sub_result;
        -- when "1110000010" => 
-- LongRes(122) <= sub_result;
        -- when "1110000011" => 
-- LongRes(121) <= sub_result;
        -- when "1110000100" => 
-- LongRes(120) <= sub_result;
        -- when "1110000101" => 
-- LongRes(119) <= sub_result;
        -- when "1110000110" => 
-- LongRes(118) <= sub_result;
        -- when "1110000111" => 
-- LongRes(117) <= sub_result;
        -- when "1110001000" => 
-- LongRes(116) <= sub_result;
        -- when "1110001001" => 
-- LongRes(115) <= sub_result;
        -- when "1110001010" => 
-- LongRes(114) <= sub_result;
        -- when "1110001011" => 
-- LongRes(113) <= sub_result;
        -- when "1110001100" => 
-- LongRes(112) <= sub_result;
        -- when "1110001101" => 
-- LongRes(111) <= sub_result;
        -- when "1110001110" => 
-- LongRes(110) <= sub_result;
        -- when "1110001111" => 
-- LongRes(109) <= sub_result;
        -- when "1110010000" => 
-- LongRes(108) <= sub_result;
        -- when "1110010001" => 
-- LongRes(107) <= sub_result;
        -- when "1110010010" => 
-- LongRes(106) <= sub_result;
        -- when "1110010011" => 
-- LongRes(105) <= sub_result;
        -- when "1110010100" => 
-- LongRes(104) <= sub_result;
        -- when "1110010101" => 
-- LongRes(103) <= sub_result;
        -- when "1110010110" => 
-- LongRes(102) <= sub_result;
        -- when "1110010111" => 
-- LongRes(101) <= sub_result;
        -- when "1110011000" => 
-- LongRes(100) <= sub_result;
        -- when "1110011001" => 
-- LongRes(99) <= sub_result;
        -- when "1110011010" => 
-- LongRes(98) <= sub_result;
        -- when "1110011011" => 
-- LongRes(97) <= sub_result;
        -- when "1110011100" => 
-- LongRes(96) <= sub_result;
        -- when "1110011101" => 
-- LongRes(95) <= sub_result;
        -- when "1110011110" => 
-- LongRes(94) <= sub_result;
        -- when "1110011111" => 
-- LongRes(93) <= sub_result;
        -- when "1110100000" => 
-- LongRes(92) <= sub_result;
        -- when "1110100001" => 
-- LongRes(91) <= sub_result;
        -- when "1110100010" => 
-- LongRes(90) <= sub_result;
        -- when "1110100011" => 
-- LongRes(89) <= sub_result;
        -- when "1110100100" => 
-- LongRes(88) <= sub_result;
        -- when "1110100101" => 
-- LongRes(87) <= sub_result;
        -- when "1110100110" => 
-- LongRes(86) <= sub_result;
        -- when "1110100111" => 
-- LongRes(85) <= sub_result;
        -- when "1110101000" => 
-- LongRes(84) <= sub_result;
        -- when "1110101001" => 
-- LongRes(83) <= sub_result;
        -- when "1110101010" => 
-- LongRes(82) <= sub_result;
        -- when "1110101011" => 
-- LongRes(81) <= sub_result;
        -- when "1110101100" => 
-- LongRes(80) <= sub_result;
        -- when "1110101101" => 
-- LongRes(79) <= sub_result;
        -- when "1110101110" => 
-- LongRes(78) <= sub_result;
        -- when "1110101111" => 
-- LongRes(77) <= sub_result;
        -- when "1110110000" => 
-- LongRes(76) <= sub_result;
        -- when "1110110001" => 
-- LongRes(75) <= sub_result;
        -- when "1110110010" => 
-- LongRes(74) <= sub_result;
        -- when "1110110011" => 
-- LongRes(73) <= sub_result;
        -- when "1110110100" => 
-- LongRes(72) <= sub_result;
        -- when "1110110101" => 
-- LongRes(71) <= sub_result;
        -- when "1110110110" => 
-- LongRes(70) <= sub_result;
        -- when "1110110111" => 
-- LongRes(69) <= sub_result;
        -- when "1110111000" => 
-- LongRes(68) <= sub_result;
        -- when "1110111001" => 
-- LongRes(67) <= sub_result;
        -- when "1110111010" => 
-- LongRes(66) <= sub_result;
        -- when "1110111011" => 
-- LongRes(65) <= sub_result;
        -- when "1110111100" => 
-- LongRes(64) <= sub_result;
        -- when "1110111101" => 
-- LongRes(63) <= sub_result;
        -- when "1110111110" => 
-- LongRes(62) <= sub_result;
        -- when "1110111111" => 
-- LongRes(61) <= sub_result;
        -- when "1111000000" => 
-- LongRes(60) <= sub_result;
        -- when "1111000001" => 
-- LongRes(59) <= sub_result;
        -- when "1111000010" => 
-- LongRes(58) <= sub_result;
        -- when "1111000011" => 
-- LongRes(57) <= sub_result;
        -- when "1111000100" => 
-- LongRes(56) <= sub_result;
        -- when "1111000101" => 
-- LongRes(55) <= sub_result;
        -- when "1111000110" => 
-- LongRes(54) <= sub_result;
        -- when "1111000111" => 
-- LongRes(53) <= sub_result;
        -- when "1111001000" => 
-- LongRes(52) <= sub_result;
        -- when "1111001001" => 
-- LongRes(51) <= sub_result;
        -- when "1111001010" => 
-- LongRes(50) <= sub_result;
        -- when "1111001011" => 
-- LongRes(49) <= sub_result;
        -- when "1111001100" => 
-- LongRes(48) <= sub_result;
        -- when "1111001101" => 
-- LongRes(47) <= sub_result;
        -- when "1111001110" => 
-- LongRes(46) <= sub_result;
        -- when "1111001111" => 
-- LongRes(45) <= sub_result;
        -- when "1111010000" => 
-- LongRes(44) <= sub_result;
        -- when "1111010001" => 
-- LongRes(43) <= sub_result;
        -- when "1111010010" => 
-- LongRes(42) <= sub_result;
        -- when "1111010011" => 
-- LongRes(41) <= sub_result;
        -- when "1111010100" => 
-- LongRes(40) <= sub_result;
        -- when "1111010101" => 
-- LongRes(39) <= sub_result;
        -- when "1111010110" => 
-- LongRes(38) <= sub_result;
        -- when "1111010111" => 
-- LongRes(37) <= sub_result;
        -- when "1111011000" => 
-- LongRes(36) <= sub_result;
        -- when "1111011001" => 
-- LongRes(35) <= sub_result;
        -- when "1111011010" => 
-- LongRes(34) <= sub_result;
        -- when "1111011011" => 
-- LongRes(33) <= sub_result;
        -- when "1111011100" => 
-- LongRes(32) <= sub_result;
        -- when "1111011101" => 
-- LongRes(31) <= sub_result;
        -- when "1111011110" => 
-- LongRes(30) <= sub_result;
        -- when "1111011111" => 
-- LongRes(29) <= sub_result;
        -- when "1111100000" => 
-- LongRes(28) <= sub_result;
        -- when "1111100001" => 
-- LongRes(27) <= sub_result;
        -- when "1111100010" => 
-- LongRes(26) <= sub_result;
        -- when "1111100011" => 
-- LongRes(25) <= sub_result;
        -- when "1111100100" => 
-- LongRes(24) <= sub_result;
        -- when "1111100101" => 
-- LongRes(23) <= sub_result;
        -- when "1111100110" => 
-- LongRes(22) <= sub_result;
        -- when "1111100111" => 
-- LongRes(21) <= sub_result;
        -- when "1111101000" => 
-- LongRes(20) <= sub_result;
        -- when "1111101001" => 
-- LongRes(19) <= sub_result;
        -- when "1111101010" => 
-- LongRes(18) <= sub_result;
        -- when "1111101011" => 
-- LongRes(17) <= sub_result;
        -- when "1111101100" => 
-- LongRes(16) <= sub_result;
        -- when "1111101101" => 
-- LongRes(15) <= sub_result;
        -- when "1111101110" => 
-- LongRes(14) <= sub_result;
        -- when "1111101111" => 
-- LongRes(13) <= sub_result;
        -- when "1111110000" => 
-- LongRes(12) <= sub_result;
        -- when "1111110001" => 
-- LongRes(11) <= sub_result;
        -- when "1111110010" => 
-- LongRes(10) <= sub_result;
        -- when "1111110011" => 
-- LongRes(9) <= sub_result;
        -- when "1111110100" => 
-- LongRes(8) <= sub_result;
        -- when "1111110101" => 
-- LongRes(7) <= sub_result;
        -- when "1111110110" => 
-- LongRes(6) <= sub_result;
        -- when "1111110111" => 
-- LongRes(5) <= sub_result;
        -- when "1111111000" => 
-- LongRes(4) <= sub_result;
        -- when "1111111001" => 
-- LongRes(3) <= sub_result;
        -- when "1111111010" => 
-- LongRes(2) <= sub_result;
        -- when "1111111011" => 
-- LongRes(1) <= sub_result;
        -- when "1111111100" => 
-- LongRes(0) <= sub_result;
         -- when others =>
     -- end case;
 -- end if;
-- end process;	
	
-- end a2;
