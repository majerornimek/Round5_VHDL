library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
use ieee.numeric_std.all;

library work;
use work.Round5_constants.all;

entity Mul_Poly_TB is
end entity; 

architecture a1 of Mul_Poly_TB is 
component Mul_Poly is 
	port (
		PolyA	: in NTRUPoly(PolyDegree downto 0);
		PolyB	: in Trinomial(PolyDegree downto 0); 
		clk		: in std_logic;
		Start	: in std_logic;
		Rst		: in std_logic;
		OpType	: in std_logic;
		Done	: out std_logic;
		LongRes	: out NTRUPoly(PolyDegree downto 0);
		ShortRes: out ShortPoly(PolyDegree downto 0)
	);
end component;
signal inA, outC : NTRUPoly(PolyDegree downto 0);
signal inB : Trinomial(PolyDegree downto  0); 
signal outS : ShortPoly(PolyDegree downto  0);
signal clk, start_tmp, rst_tmp, op_tmp, done_tmp : std_logic;
constant CLK_PERIOD : time := 10 ps;
type input_array is array(PolyDegree downto 0) of integer;

begin

 clk_process :process
   begin
        clk <= '0';
        wait for CLK_PERIOD/2;  --for half of clock period clk stays at '0'.
        clk <= '1';
        wait for CLK_PERIOD/2;  --for next half of clock period clk stays at '1'.
   end process;
   
   uut: Mul_Poly port map(
    	PolyA	=> inA,
		PolyB	=> inB,
		clk		=> clk,
		Start	=> start_tmp,
		Rst		=> rst_tmp,
		OpType	=> op_tmp,
		Done	=> done_tmp,
		LongRes	=> outC,
		ShortRes=> outS
   );
   
process
	
	procedure check_poly_mul( 	constant PolyA	: in input_array; -- v1
								constant PolyB 	: in input_array; -- v2
								constant typ	: in std_logic; -- norm of v1
								constant res_ex	: in input_array) is
		variable res: input_array;
	begin
		GG: for i in PolyDegree downto 0 loop
			inA(i) <= std_logic_vector(to_signed(PolyA(i), LongModLen-1));
			inB(i) <= std_logic_vector(to_signed(PolyB(i), 2));
		end loop GG; 
		
		wait for CLK_PERIOD;
		rst_tmp <= '1';
		op_tmp <= typ;
		wait for CLK_PERIOD;
		rst_tmp <= '0';
		start_tmp <= '1';
		wait for CLK_PERIOD*1400;
		start_tmp <= '0';
		wait for CLK_PERIOD;
		
--		RR: for i in NUM_OF_ELEMENTS-1 downto 0 loop
--			res(i) = to_integer(signed(outC(i)));
--		end loop RR;
--		assert res = res_ex
--		report 	"Unexpected result: " --&
----				"IN1 = " & integer'image(in1) & "; " &
----				"IN2 = " & integer'image(in2) & "; " &
----				"MUL = " & integer'image(res) & "; " &
----				"MUL_expected = " & integer'image(res_ex)
--		severity error;
	end procedure check_poly_mul;
	
	
begin
	
    check_poly_mul((784,2028,1705,574,571,1226,1324,236,642,1876,105,1158,388,1119,1563,204,1977,1595,1048,1785,1845,1345,1894,1990,1591,1753,1276,1568,104,1220,651,511,38,1343,701,1517,402,1727,291,438,381,101,506,35,120,1370,806,362,953,1959,805,606,457,13,1037,1904,614,1745,703,2027,813,1634,2017,917,1269,910,717,497,1325,2017,1869,266,992,1904,204,1208,1363,801,799,1535,965,1104,253,1493,1360,122,1850,1903,1775,1021,972,1961,1545,1390,255,595,1105,1037,937,689,802,1039,1930,1728,134,1894,1650,1230,294,1382,651,1966,1544,459,947,1983,491,648,1363,2040,279,50,880,700,301,816,319,934,1204,263,1196,1348,1395,1059,1238,942,69,1105,319,266,1794,1591,1264,439,1462,1244,1812,1404,1920,153,653,61,299,411,1528,404,745,12,894,1573,961,1716,1725,863,1623,906,1992,188,1297,1113,1829,573,949,627,1733,1247,739,777,1926,1765,1630,991,1574,1567,5,1955,693,19,1594,424,509,1947,1761,1201,263,1565,119,1736,1755,349,784,447,1495,455,400,1636,1731,702,1610,1959,964,1396,1673,1970,443,303,1369,959,574,809,719,1659,771,1709,1756,1421,1992,672,1648,792,189,1181,275,466,1171,153,1101,354,969,348,1217,1452,2043,734,1930,1056,1042,1218,218,1313,362,43,945,825,332,1334,707,23,283,904,779,1830,404,1772,1677,1933,574,352,98,762,1384,1433,1717,1455,512,528,1423,435,693,856,116,659,381,129,308,1242,373,86,735,1841,995,1278,1563,669,485,147,1043,2026,1648,1615,934,186,616,2008,1698,314,963,699,148,1271,538,1037,968,947,606,822,1944,1053,1498,1765,1974,1310,352,790,411,1743,1529,142,1514,565,1190,450,164,487,1135,733,15,626,545,1039,828,678,1350,727,791,1909,1314,660,1223,1209,1097,448,1467,603,1352,1836,1854,360,1668,212,1403,1227,461,411,2031,408,1115,38,554,874,1916,1858,2033,1777,1754,1542,1220,1704,1645,1040,366,1279,864,15,932,570,796,692,1342,99,877,713,9,1474,267,501,175,1612,769,1877,831,870,888,1656,231,129,987,560,1611,1828,113,621,1370,786,272,677,718,419,1141,1029,622,549,277,1003,1500,1876,487,320,1429,951,365,1899,138,1162,1625,863,1848,735,15,187,1288,317,1019,663,1591,1987,597,1654,296,1519,1277,1099,954,1891,1904,935,910,2045,149,1735,679,507,1125,221,75,1016,1541,656,750,1717,1585,212,1035,1965,328,1263,1054,1634,968,1512,1269,1334,2045,1783,1306,268,971,1649,126,572,1118,186,1574,1623,1048,1451,289,1785,1563,999,1053,1007,547,586,291,1690,211,255,409,647,325,1951,676,995,59,1841,1239,1026,1509,141,224,772,520,376,125,1039,1598,1141,159,1931,79,1709,1349,475,132,1109,705,916,1261,1331,316,22,904,1670,955,1764,276,285,385,1525,457,823,1392,478,1557,1382,23,1165,500,1272,564,393,442,138,1891,1513,1405,1982,175,895,701,1022,1828,981,50,846,489,1668,885,477,175,991,1089,728,640,724,247,950,1930,644,2016,1174,1857,1061,239,1819,1809,1529,1391,1062,523,1469,1849,154,291,1939,1672,912,1682,840,1730,89,300,1405,1288,374,1021,985,0),
    (0,0,0,0,0,0,0,-1,0,0,0,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,1,0,0,1,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,1,-1,0,0,0,-1,0,0,-1,0,0,0,0,0,0,0,1,0,1,0,0,1,0,0,0,0,0,0,0,-1,1,1,0,0,0,0,0,1,0,0,0,0,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,0,0,0,0,0,0,-1,0,0,0,0,0,0,1,0,0,1,0,0,0,1,0,0,0,0,0,0,0,0,0,0,-1,1,-1,0,0,0,0,0,1,0,0,-1,0,0,0,0,0,0,0,0,0,1,-1,0,1,0,0,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,0,0,0,0,-1,0,-1,0,0,0,1,-1,0,0,0,0,0,0,0,0,-1,0,-1,0,0,0,0,0,-1,0,0,0,0,0,-1,0,0,1,0,0,0,0,0,0,0,0,0,0,-1,0,1,1,0,0,0,0,0,0,0,0,0,0,-1,-1,1,1,0,0,0,0,0,0,1,0,0,-1,-1,0,0,0,0,0,0,1,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,-1,0,0,0,-1,0,0,1,0,0,0,0,1,0,0,0,0,0,0,0,0,0,-1,0,1,0,0,0,0,0,0,0,1,0,0,0,-1,1,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,0,0,1,1,0,0,0,0,0,0,0,-1,0,0,1,1,0,0,0,0,0,0,0,1,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,0,0,0,0,0,0,0,0,0,0,-1,0,0,-1,0,0,-1,0,0,0,0,-1,1,-1,0,0,0,0,0,0,0,-1,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,1,0,0,0,0,0,0,0,0,0,0,-1,0,-1,-1,0,1,0,0,0,0,0,0,0,0,0,0,1,0,1,1,-1,-1,0,0,0,0,0,0,-1,0,0,0,0,0,0,0,0,1,0,0,0,0,-1,0,0,0,0),
   '1',
	(0,589, 1400, 1227, 1545, 1045, 1921, 109, 1569, 108, 1754, 1556, 14, 1409, 237, 1106, 1922, 1259, 1966, 583, 747, 510, 1545, 1994, 35, 1613, 1439, 1064, 1147, 730, 1932, 1819, 1580, 1517, 324, 1459, 161, 600, 711, 530, 503, 784, 912, 14, 562, 739, 1649, 609, 346, 1695, 405, 928, 2034, 1988, 1541, 1761, 156, 833, 1503, 112, 1486, 854, 588, 871, 616, 127, 1865, 1837, 2034, 961, 1861, 193, 521, 1206, 471, 788, 517, 1436, 603, 1692, 1558, 1329, 1576, 1641, 2003, 1193, 1339, 1665, 1553, 58, 2003, 1981, 256, 267, 1760, 690, 1879, 1954, 1905, 1516, 1834, 284, 218, 421, 1, 1030, 416, 97, 121, 1175, 1816, 1663, 1754, 249, 1462, 1305, 2029, 1977, 1497, 1713, 669, 642, 593, 1462, 1085, 1306, 1498, 547, 1385, 1961, 1113, 910, 1786, 432, 564, 825, 658, 763, 1529, 460, 901, 1815, 1810, 956, 853, 1824, 361, 558, 1973, 1948, 1687, 1673, 45, 1548, 847, 1220, 1873, 578, 482, 1035, 760, 1383, 1224, 1907, 1287, 918, 897, 1454, 573, 2017, 1548, 317, 641, 1019, 525, 1286, 48, 1132, 1227, 1907, 75, 1180, 366, 1871, 1568, 1658, 718, 110, 107, 1256, 536, 1788, 360, 792, 257, 928, 1872, 831, 42, 610, 1724, 286, 908, 1266, 326, 1827, 1444, 1927, 889, 1405, 1270, 1757, 1617, 296, 1753, 1628, 1144, 1543, 1529, 1209, 808, 1399, 443, 1564, 1381, 323, 1277, 91, 1269, 1553, 453, 1466, 1443, 443, 2042, 1923, 1559, 834, 1897, 281, 251, 312, 455, 1510, 563, 260, 1714, 1337, 348, 1691, 1624, 1601, 1027, 1552, 914, 746, 630, 1287, 66, 467, 1932, 1053, 513, 310, 1164, 612, 93, 488, 1945, 40, 882, 506, 221, 1831, 547, 1158, 1398, 1147, 1781, 1051, 1608, 1925, 1870, 1404, 922, 1413, 2, 876, 1252, 591, 301, 818, 995, 1659, 854, 740, 1391, 1225, 1420, 1842, 714, 1478, 1154, 1619, 286, 2029, 273, 516, 1754, 1980, 1636, 13, 243, 43, 1873, 151, 1659, 228, 437, 351, 463, 1826, 379, 881, 1155, 1658, 1646, 576, 1771, 1410, 447, 1674, 480, 1423, 35, 1916, 746, 1799, 721, 138, 1536, 280, 1955, 853, 663, 47, 1734, 653, 801, 561, 1518, 1401, 587, 518, 41, 214, 239, 1932, 28, 1781, 1377, 1251, 260, 958, 64, 380, 2015, 163, 171, 1351, 15, 129, 850, 683, 252, 1623, 100, 1245, 443, 1658, 874, 1547, 1312, 1437, 1730, 510, 635, 1391, 230, 1197, 1130, 740, 1097, 1644, 1145, 1625, 1410, 525, 1245, 1124, 1523, 1823, 1642, 1356, 1708, 133, 1811, 723, 1565, 1241, 928, 185, 1168, 2041, 259, 653, 113, 817, 1875, 1490, 1005, 622, 2032, 919, 734, 133, 1998, 93, 1910, 983, 484, 1445, 276, 226, 1090, 1161, 409, 1928, 1276, 1580, 841, 1494, 716, 1613, 1838, 1349, 518, 1755, 2014, 692, 1783, 668, 1282, 1772, 1008, 1343, 358, 1249, 1906, 108, 285, 1043, 1522, 1167, 1901, 15, 1542, 1866, 1998, 233, 1055, 959, 993, 1301, 1421, 2002, 962, 662, 731, 1299, 728, 384, 1510, 130, 503, 1031, 346, 1022, 1404, 152, 1257, 158, 1734, 1840, 671, 833, 733, 1232, 1035, 139, 680, 1494, 1830, 642, 567, 1704, 1019, 1370, 1874, 495, 1122, 1380, 237, 1851, 332, 336, 1853, 1470, 1383, 1242, 279, 1200, 1431, 864, 367, 973, 297, 269, 1708, 852, 880, 1965, 663, 228, 40, 837, 1359, 446, 306, 1262, 1573, 784, 186, 1302, 344, 1185, 342, 388, 892, 1887, 1216, 1602, 1498, 79, 347, 1643, 1162, 929, 434, 1914, 674, 903, 1709, 1931, 1904, 283, 1734, 367, 1991, 504, 667, 1135, 1951, 1873, 29, 1872, 1061, 890, 436, 2028, 995, 459, 602, 674, 939, 1509, 830, 1724, 42, 1224, 1003, 1305, 342, 1355, 804, 1099, 52, 677, 181, 1629, 2017, 1633, 339, 1316, 352, 247, 9, 1072, 1314, 1512, 1077, 87, 220, 1067, 124, 1614, 1291, 776, 1398)
   );
end process;   
   
end a1;