library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
use ieee.numeric_std.all;
--use ieee.std_logic_arith.all;

library work;
use work.Round5_constants.all;

entity Round5_enc_arith_TB is	
end entity;

architecture a1 of Round5_enc_arith_TB is

component Round5_enc_arith is	
	port (
		PolyA			: in q_bitsPoly(PolyDegree-1 downto 0);  --W enc: A
		PolyB			: in p_bitsPoly(PolyDegree downto 0);	--W enc: polyB,   W dec: polyU
		PolyR			: in Trinomial(PolyDegree-1 downto 0); --W enc: poly R   W dec: polyS
		Message		: in std_logic_vector(MessageLen-1 downto 0);
		
		clk			: in std_logic;
		Start			: in std_logic;
		Reset			: in std_logic;
		Operation	: in std_logic;  -- 1 enc, 0 dec
		
		FirstPart	: out p_bitsPoly(PolyDegree-1 downto 0);
		SecondPart	: out t_bitsPoly(PolyDegree-1 downto 0)
	);
end component;

signal clk : std_logic;

constant CLK_PERIOD : time := 10 ps;
signal PolyA_tmp, Result_tmp : q_bitsPoly(PolyDegree-1 downto 0);
signal PolyB_tmp : p_bitsPoly(PolyDegree downto 0);
signal PolyR_tmp : Trinomial(PolyDegree-1 downto 0);
signal Message_tmp : std_logic_vector(MessageLen-1 downto 0);


signal short_Res : p_bitsPoly(PolyDegree downto 0);
signal start_tmp, reset_tmp, op_tmp : std_logic;
type input_array is array(PolyDegree-1 downto 0) of integer;
type input_array2 is array(PolyDegree downto 0) of integer;
signal first_tmp :p_bitsPoly(PolyDegree-1 downto 0);
signal second_tmp : t_bitsPoly(PolyDegree-1 downto 0);
signal b1,b2,b3 : input_array;
--
--constant c1 : input_array := 1203, 1807, 1535, 215, 11, 1536, 1011, 1996, 68, 622, 926, 1641, 744, 1729, 74, 1004, 276, 239, 1713, 1601, 1075, 1175, 417, 688, 479, 1892, 1478, 121, 1162, 94, 831, 1159, 1515, 1499, 1861, 1763, 1543, 1992, 1618, 1404, 1619, 1874, 483, 1238, 170, 1514, 1199, 2006, 1187, 66, 313, 452, 1049, 789, 1964, 1866, 1788, 137, 1571, 721, 736, 996, 171, 1728, 1219, 1837, 1400, 1027, 199, 786, 360, 1580, 1174, 914, 273, 92, 111, 1984, 1087, 781, 452, 1423, 202, 295, 1515, 391, 1712, 1112, 1902, 1814, 399, 455, 385, 1715, 651, 987, 1723, 1545, 1575, 1351, 538, 109, 859, 721, 1821, 571, 1261, 1846, 1622, 613, 1892, 1198, 1952, 218, 357, 64, 1824, 325, 573, 219, 1481, 919, 899, 693, 1636, 1966, 140, 302, 219, 232, 1083, 582, 577, 964, 1680, 1941, 842, 483, 850, 1090, 1192, 758, 1767, 59, 459, 1218, 1760, 1800, 608, 1354, 3, 1903, 329, 1480, 1618, 1764, 1597, 1279, 188, 1908, 1896, 937, 1370, 1413, 1669, 1467, 167, 1480, 1185, 228, 1051, 90, 1393, 466, 1467, 509, 271, 1982, 771, 2046, 2030, 795, 653, 1570, 128, 1808, 1594, 658, 1752, 1256, 1813, 1172, 240, 1267, 1457, 1006, 1096, 38, 112, 1469, 960, 1305, 10, 674, 1562, 1573, 1344, 1472, 1111, 1280, 1060, 668, 1049, 901, 733, 1819, 1944, 32, 595, 515, 1692, 47, 942, 1735, 463, 951, 1350, 1253, 1073, 1019, 1701, 1564, 1237, 1269, 1564, 27, 1147, 870, 919, 113, 903, 1422, 287, 1718, 1879, 1335, 57, 1237, 516, 340, 1223, 1697, 205, 1278, 1474, 1407, 1924, 967, 1515, 1999, 1805, 1596, 51, 310, 1369, 322, 595, 215, 594, 716, 1447, 1505, 176, 1302, 315, 2004, 1895, 385, 470, 1668, 368, 534, 1290, 1761, 174, 63, 1177, 415, 1641, 1650, 356, 1090, 700, 1612, 1662, 937, 577, 1014, 1689, 480, 1449, 1229, 625, 2044, 2022, 1820, 908, 1233, 1148, 804, 1950, 1950, 164, 216, 191, 1569, 78, 1885, 1429, 568, 836, 2043, 1121, 1579, 1023, 2036, 596, 1441, 1643, 1267, 1830, 1145, 846, 1976, 1184, 1515, 1072, 1690, 1533, 1598, 330, 281, 1024, 1729, 1798, 1080, 1736, 861, 1423, 1812, 795, 1015, 1296, 552, 1069, 921, 64, 2026, 799, 409, 521, 1917, 348, 841, 1344, 1142, 1523, 822, 520, 300, 877, 397, 1131, 1816, 1483, 1587, 1097, 1391, 1623, 943, 628, 986, 418, 106, 1689, 1949, 1629, 222, 1201, 1133, 616, 1321, 970, 1555, 457, 532, 1500, 1329, 471, 263, 168, 1079, 648, 695, 647, 1602, 1834, 140, 1148, 937, 1750, 1839, 1534, 975, 683, 1539, 1945, 633, 1160, 297, 1944, 1844, 1802, 532, 1630, 1334, 1040, 196, 456, 569, 391, 1229, 749, 1138, 288, 1630, 565, 1223, 1061, 833, 1573, 1430, 127, 1761, 1249, 687, 1070, 82, 1145, 1272, 1552, 1023, 214, 253, 376, 1169, 1855, 81, 578, 1461, 914, 1717, 1889, 5, 1755, 1570, 1729, 324, 643, 1671, 866, 1429, 886, 1568, 1828, 1399, 1564, 397, 1612, 972, 831, 300, 830, 1317, 31, 1537, 19, 1762, 1747, 32, 1413, 1990, 458, 852, 453, 56, 1194, 1436, 112, 799, 1692, 187, 1824, 20, 923, 1818, 1813, 814, 1282, 1409, 493, 937, 1260, 1041, 4, 1848, 169, 662, 48, 1972, 1380, 380, 1004, 1841, 1175, 1401, 1254, 196, 1797, 346, 552, 2013, 963, 81, 1684, 1702, 1250, 358, 1588, 495, 1620, 1306, 1150, 223, 1773, 1109, 825, 1896, 135, 1424, 1257, 1911, 177, 1860, 1392, 663, 1921, 6, 1019, 1239, 1925, 1179, 362, 1215, 1115, 1288, 1128, 900, 334, 1406, 1880, 406, 872, 1943, 1256, 1425, 1096, 88, 1586, 26, 1087, 835, 1943, 1784, 1387, 1225, 521, 675, 681, 1549, 143, 1475, 1077, 1553, 894, 798, 1349, 1885, 1162, 1911, 120, 1110, 1718, 635, 942, 230, 1152, 154, 1215, 1430, 1521, 780, 1833, 1161, 47, 977, 714, 306),		(62, 119, 242, 38, 67, 246, 55, 252, 233, 46, 101, 25, 165, 21, 141, 246, 126, 85, 8, 35, 78, 148, 28, 178, 247, 154, 230, 5, 96, 196, 242, 175, 234, 12, 212, 114, 56, 73, 40, 60, 2, 24, 187, 123, 176, 233, 143, 13, 142, 45, 179, 82, 177, 243, 120, 104, 252, 229, 91, 114, 148, 249, 129, 59, 162, 9, 127, 49, 96, 197, 181, 203, 118, 11, 16, 164, 65, 1, 89, 110, 112, 125, 12, 101, 32, 117, 76, 122, 231, 100, 146, 235, 84, 167, 78, 140, 166, 137, 214, 253, 3, 240, 105, 246, 102, 55, 252, 24, 51, 246, 25, 113, 140, 130, 107, 208, 246, 70, 147, 222, 52, 12, 214, 217, 170, 1, 175, 210, 226, 161, 178, 143, 51, 240, 226, 16, 213, 91, 237, 232, 84, 8, 20, 219, 247, 78, 241, 218, 216, 208, 211, 121, 167, 39, 165, 253, 151, 119, 131, 170, 166, 222, 56, 204, 200, 138, 184, 23, 72, 91, 0, 132, 42, 117, 211, 155, 71, 240, 33, 117, 146, 178, 169, 253, 119, 121, 125, 224, 29, 70, 159, 81, 136, 29, 169, 145, 24, 87, 161, 60, 119, 127, 155, 250, 237, 128, 213, 144, 54, 126, 65, 151, 251, 47, 221, 77, 237, 19, 134, 44, 228, 150, 176, 181, 133, 50, 242, 159, 119, 106, 159, 81, 21, 43, 247, 247, 137, 41, 72, 246, 150, 139, 124, 16, 165, 97, 176, 62, 65, 217, 194, 84, 158, 255, 185, 113, 241, 29, 248, 33, 55, 53, 245, 160, 170, 178, 187, 40, 125, 54, 206, 34, 94, 101, 108, 93, 136, 97, 100, 79, 220, 90, 255, 232, 254, 29, 159, 58, 25, 4, 202, 166, 237, 246, 147, 229, 210, 84, 126, 175, 136, 42, 224, 154, 225, 32, 52, 198, 126, 69, 221, 142, 167, 226, 15, 184, 209, 185, 95, 20, 115, 22, 65, 140, 173, 89, 42, 31, 42, 67, 107, 182, 217, 211, 90, 5, 19, 15, 192, 165, 246, 90, 155, 5, 212, 157, 103, 36, 232, 202, 145, 185, 141, 177, 247, 30, 226, 80, 57, 63, 9, 116, 27, 113, 251, 33, 171, 201, 103, 84, 80, 144, 117, 104, 138, 6, 188, 226, 156, 201, 43, 130, 109, 135, 139, 225, 169, 7, 160, 242, 6, 185, 129, 114, 37, 205, 131, 6, 89, 42, 92, 100, 221, 150, 81, 225, 66, 201, 23, 245, 43, 69, 46, 89, 248, 35, 38, 171, 63, 12, 173, 135, 128, 30, 41, 107, 92, 231, 183, 11, 254, 9, 80, 69, 120, 92, 165, 152, 4, 158, 54, 233, 56, 64, 86, 165, 160, 93, 178, 154, 83, 101, 53, 37, 66, 240, 195, 235, 132, 183, 139, 121, 181, 213, 63, 88, 93, 42, 234, 136, 198, 132, 136, 175, 211, 241, 252, 36, 143, 143, 209, 132, 178, 215, 166, 177, 80, 197, 176, 25, 225, 231, 179, 249, 168, 155, 93, 250, 34, 156, 219, 255, 163, 24, 128, 234, 206, 232, 232, 8, 146, 242, 123, 176, 48, 24, 169, 171, 238, 197, 211, 34, 39, 177, 126, 154, 142, 170, 70, 176, 237, 15, 250, 67, 240, 17, 187, 15, 184, 177, 7, 111, 111, 186, 217, 101, 243, 131, 121, 152, 162, 156, 59, 98, 237, 251, 25, 146, 54, 47, 43, 237, 44, 15, 14, 73, 253, 39, 201, 210, 36, 19, 183, 32, 33, 3, 141, 105, 233, 174, 33, 168, 159, 235, 132, 3, 63, 242, 193, 126, 208, 4, 241, 85, 210, 72, 230, 95, 60, 224, 109, 237, 88, 115, 135, 59, 78, 90, 226, 146, 181, 0, 45, 78, 45, 123, 15, 137;
--constant c2 : input_array := (165, 57, 101, 115, 149, 111, 165, 88, 187, 42, 121, 5, 218, 100, 241, 200, 201, 181, 226, 249, 149, 68, 118, 182, 40, 120, 36, 110, 62, 12, 63, 142, 109, 194, 25, 28, 94, 1, 90, 167, 117, 40, 88, 53, 116, 155, 78, 120, 136, 183, 103, 68, 141, 192, 18, 11, 187, 167, 147, 58, 80, 248, 125, 236, 176, 163, 238, 95, 30, 3, 82, 248, 21, 203, 144, 240, 167, 197, 63, 182, 209, 50, 162, 3, 241, 113, 193, 196, 198, 217, 32, 20, 224, 2, 90, 236, 254, 231, 19, 105, 84, 94, 226, 210, 251, 56, 124, 193, 225, 220, 160, 249, 13, 159, 154, 119, 84, 101, 212, 107, 22, 236, 210, 101, 43, 167, 89, 246, 185, 132, 29, 13, 99, 203, 93, 158, 122, 220, 4, 251, 138, 104, 229, 131, 32, 212, 26, 250, 189, 193, 194, 138, 246, 13, 6, 35, 128, 55, 94, 22, 171, 209, 133, 58, 208, 72, 114, 84, 238, 43, 207, 156, 154, 87, 34, 29, 165, 39, 128, 103, 143, 101, 194, 13, 64, 192, 213, 94, 149, 253, 99, 79, 8, 29, 150, 247, 135, 205, 121, 244, 99, 63, 36, 118, 2, 133, 217, 69, 72, 122, 59, 99, 39, 241, 136, 214, 108, 138, 179, 238, 185, 195, 142, 2, 165, 128, 165, 202, 227, 251, 136, 184, 98, 206, 228, 157, 69, 59, 178, 147, 195, 72, 147, 9, 207, 85, 218, 104, 221, 19, 172, 90, 218, 192, 71, 199, 135, 206, 209, 92, 141, 150, 182, 225, 161, 7, 154, 92, 173, 3, 37, 143, 75, 150, 145, 90, 219, 58, 192, 92, 175, 159, 227, 9, 233, 155, 243, 207, 151, 197, 72, 78, 125, 143, 255, 71, 252, 197, 36, 198, 209, 34, 129, 228, 72, 206, 19, 95, 115, 15, 20, 0, 85, 104, 10, 61, 53, 62, 63, 60, 122, 243, 122, 144, 47, 139, 80, 251, 72, 96, 33, 13, 116, 172, 70, 81, 113, 243, 118, 243, 7, 193, 186, 56, 124, 237, 12, 206, 6, 159, 13, 58, 240, 227, 91, 191, 201, 254, 75, 192, 135, 244, 147, 101, 250, 134, 153, 75, 236, 95, 113, 27, 133, 81, 222, 108, 7, 196, 190, 23, 163, 182, 185, 30, 102, 228, 170, 36, 28, 90, 161, 30, 4, 222, 215, 181, 30, 225, 57, 118, 93, 212, 47, 180, 7, 156, 98, 81, 222, 247, 218, 55, 90, 67, 34, 188, 224, 56, 234, 68, 158, 39, 242, 239, 8, 124, 248, 59, 190, 55, 147, 26, 244, 4, 141, 202, 139, 144, 169, 243, 101, 102, 95, 170, 201, 105, 17, 50, 176, 142, 61, 175, 83, 2, 111, 165, 93, 76, 29, 123, 136, 15, 187, 243, 55, 71, 238, 28, 46, 13, 91, 61, 162, 34, 119, 59, 238, 205, 244, 92, 159, 196, 117, 180, 32, 177, 122, 19, 24, 228, 137, 128, 173, 173, 20, 0, 250, 39, 214, 146, 64, 76, 43, 48, 85, 207, 37, 119, 55, 208, 171, 82, 5, 231, 50, 240, 129, 246, 208, 152, 96, 12, 96, 180, 61, 248, 194, 62, 231, 147, 40, 247, 201, 252, 46, 73, 115, 106, 121, 232, 77, 22, 8, 115, 61, 229, 216, 253, 246, 123, 170, 24, 252, 168, 107, 201, 188, 25, 246, 78, 218, 218, 206, 0, 174, 115, 139, 239, 85, 198, 136, 1, 65, 191, 59, 68, 188, 58, 95, 247, 226, 162, 169, 116, 172, 100, 102, 142, 166, 90, 33, 48, 208, 1, 236, 64, 162, 131, 75, 137, 147, 214, 110, 147, 149, 101, 71, 249, 137, 135, 108, 113, 74, 195, 50, 105, 240, 227);
--constant c3 : input_array := (0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, 1, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, -1, 0, 0, -1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0);

begin

	clk_process :process
   begin
        clk <= '0';
        wait for CLK_PERIOD/2;  --for half of clock period clk stays at '0'.
        clk <= '1';
        wait for CLK_PERIOD/2;  --for next half of clock period clk stays at '1'.
   end process;


	uut: Round5_enc_arith port map(
		PolyA			=> PolyA_tmp,
		PolyB			=> PolyB_tmp,
		PolyR			=> PolyR_tmp,
		Message		=> Message_tmp,
		
		clk			=> clk,
		Start			=> Start_tmp,
		Reset			=> Reset_tmp,
		Operation	=> op_tmp,
		
		FirstPart	=> first_tmp,
		SecondPart => Second_tmp
	);
	
	
	
	
	
	
process

		procedure check_enc( 	constant inV1	: in input_array; -- v1
										constant inV2	: in input_array2;
										constant inV3	: in input_array;--;
										constant inV4	: in std_logic_vector(MessageLen-1 downto 0)
									) is
									
		variable res: input_array;
		
		begin
			GG: for i in PolyDegree-1 downto 0 loop
				PolyA_tmp(i) <= std_logic_vector(to_unsigned(inV1(i), q_bits));
				PolyB_tmp(i) <= std_logic_vector(to_unsigned(inV2(i), p_bits));
				PolyR_tmp(i) <= std_logic_vector(to_signed(inV3(i), 2));
				
			end loop GG;
				PolyB_tmp(PolyDegree) <= std_logic_vector(to_unsigned(inV2(PolyDegree), p_bits));
			
				Message_tmp <= inV4;--"00111100110011001110010111100001101100100001011001101001110110101100101001011111010000111000101111011000011101011111111010000100";
				
			wait for CLK_PERIOD;
			start_tmp <= '1';
			op_tmp <= '1';
			wait for 5*CLK_PERIOD*(PolyDegree+5);
			start_tmp <= '0';
			wait for  CLK_PERIOD;
			RR: for i in PolyDegree-1 downto 0 loop
				res(i) := to_integer(unsigned(Result_tmp(i)));

			end loop RR;
			assert res /= inV1
			report 	"Unexpected result: " --&
	--				"IN1 = " & integer'image(in1) & "; " &
	--				"IN2 = " & integer'image(in2) & "; " &
	--				"MUL = " & integer'image(res) & "; " &
	--				"MUL_expected = " & integer'image(res_ex)
			severity error;
		end procedure check_enc;
        
        
        procedure check_dec( 	        constant inV1	: in input_array; --  U, short Poly, B
										constant inV2	: in input_array2;
										constant inV3	: in input_array;--;
										constant inV4	: in std_logic_vector(MessageLen-1 downto 0)
									) is
									
		variable res: input_array;
		
		begin
			GG: for i in PolyDegree-1 downto 0 loop
				PolyB_tmp(i) <= std_logic_vector(to_unsigned(inV1(i), ShortModLen-1));
				PolyR_tmp(i) <= std_logic_vector(to_signed(inV3(i), 2));
				
			end loop GG;
				PolyB_tmp(PolyDegree) <= std_logic_vector(to_unsigned(inV2(PolyDegree), ShortModLen-1));
			
				Message_tmp <= inV4;--"00111100110011001110010111100001101100100001011001101001110110101100101001011111010000111000101111011000011101011111111010000100";
				
			wait for CLK_PERIOD;
			start_tmp <= '1';
			op_tmp <= '0';
			wait for 5*CLK_PERIOD*(PolyDegree+5);
			start_tmp <= '0';
			wait for  CLK_PERIOD;
			RR: for i in PolyDegree-1 downto 0 loop
				res(i) := to_integer(unsigned(Result_tmp(i)));

			end loop RR;
			assert res /= inV1
			report 	"Unexpected result: " --&
	--				"IN1 = " & integer'image(in1) & "; " &
	--				"IN2 = " & integer'image(in2) & "; " &
	--				"MUL = " & integer'image(res) & "; " &
	--				"MUL_expected = " & integer'image(res_ex)
			severity error;
		end procedure check_dec;
        
	
	begin
		wait for CLK_PERIOD;
		start_tmp <=	'0';

		check_enc(
		(1203, 1807, 1535, 215, 11, 1536, 1011, 1996, 68, 622, 926, 1641, 744, 1729, 74, 1004, 276, 239, 1713, 1601, 1075, 1175, 417, 688, 479, 1892, 1478, 121, 1162, 94, 831, 1159, 1515, 1499, 1861, 1763, 1543, 1992, 1618, 1404, 1619, 1874, 483, 1238, 170, 1514, 1199, 2006, 1187, 66, 313, 452, 1049, 789, 1964, 1866, 1788, 137, 1571, 721, 736, 996, 171, 1728, 1219, 1837, 1400, 1027, 199, 786, 360, 1580, 1174, 914, 273, 92, 111, 1984, 1087, 781, 452, 1423, 202, 295, 1515, 391, 1712, 1112, 1902, 1814, 399, 455, 385, 1715, 651, 987, 1723, 1545, 1575, 1351, 538, 109, 859, 721, 1821, 571, 1261, 1846, 1622, 613, 1892, 1198, 1952, 218, 357, 64, 1824, 325, 573, 219, 1481, 919, 899, 693, 1636, 1966, 140, 302, 219, 232, 1083, 582, 577, 964, 1680, 1941, 842, 483, 850, 1090, 1192, 758, 1767, 59, 459, 1218, 1760, 1800, 608, 1354, 3, 1903, 329, 1480, 1618, 1764, 1597, 1279, 188, 1908, 1896, 937, 1370, 1413, 1669, 1467, 167, 1480, 1185, 228, 1051, 90, 1393, 466, 1467, 509, 271, 1982, 771, 2046, 2030, 795, 653, 1570, 128, 1808, 1594, 658, 1752, 1256, 1813, 1172, 240, 1267, 1457, 1006, 1096, 38, 112, 1469, 960, 1305, 10, 674, 1562, 1573, 1344, 1472, 1111, 1280, 1060, 668, 1049, 901, 733, 1819, 1944, 32, 595, 515, 1692, 47, 942, 1735, 463, 951, 1350, 1253, 1073, 1019, 1701, 1564, 1237, 1269, 1564, 27, 1147, 870, 919, 113, 903, 1422, 287, 1718, 1879, 1335, 57, 1237, 516, 340, 1223, 1697, 205, 1278, 1474, 1407, 1924, 967, 1515, 1999, 1805, 1596, 51, 310, 1369, 322, 595, 215, 594, 716, 1447, 1505, 176, 1302, 315, 2004, 1895, 385, 470, 1668, 368, 534, 1290, 1761, 174, 63, 1177, 415, 1641, 1650, 356, 1090, 700, 1612, 1662, 937, 577, 1014, 1689, 480, 1449, 1229, 625, 2044, 2022, 1820, 908, 1233, 1148, 804, 1950, 1950, 164, 216, 191, 1569, 78, 1885, 1429, 568, 836, 2043, 1121, 1579, 1023, 2036, 596, 1441, 1643, 1267, 1830, 1145, 846, 1976, 1184, 1515, 1072, 1690, 1533, 1598, 330, 281, 1024, 1729, 1798, 1080, 1736, 861, 1423, 1812, 795, 1015, 1296, 552, 1069, 921, 64, 2026, 799, 409, 521, 1917, 348, 841, 1344, 1142, 1523, 822, 520, 300, 877, 397, 1131, 1816, 1483, 1587, 1097, 1391, 1623, 943, 628, 986, 418, 106, 1689, 1949, 1629, 222, 1201, 1133, 616, 1321, 970, 1555, 457, 532, 1500, 1329, 471, 263, 168, 1079, 648, 695, 647, 1602, 1834, 140, 1148, 937, 1750, 1839, 1534, 975, 683, 1539, 1945, 633, 1160, 297, 1944, 1844, 1802, 532, 1630, 1334, 1040, 196, 456, 569, 391, 1229, 749, 1138, 288, 1630, 565, 1223, 1061, 833, 1573, 1430, 127, 1761, 1249, 687, 1070, 82, 1145, 1272, 1552, 1023, 214, 253, 376, 1169, 1855, 81, 578, 1461, 914, 1717, 1889, 5, 1755, 1570, 1729, 324, 643, 1671, 866, 1429, 886, 1568, 1828, 1399, 1564, 397, 1612, 972, 831, 300, 830, 1317, 31, 1537, 19, 1762, 1747, 32, 1413, 1990, 458, 852, 453, 56, 1194, 1436, 112, 799, 1692, 187, 1824, 20, 923, 1818, 1813, 814, 1282, 1409, 493, 937, 1260, 1041, 4, 1848, 169, 662, 48, 1972, 1380, 380, 1004, 1841, 1175, 1401, 1254, 196, 1797, 346, 552, 2013, 963, 81, 1684, 1702, 1250, 358, 1588, 495, 1620, 1306, 1150, 223, 1773, 1109, 825, 1896, 135, 1424, 1257, 1911, 177, 1860, 1392, 663, 1921, 6, 1019, 1239, 1925, 1179, 362, 1215, 1115, 1288, 1128, 900, 334, 1406, 1880, 406, 872, 1943, 1256, 1425, 1096, 88, 1586, 26, 1087, 835, 1943, 1784, 1387, 1225, 521, 675, 681, 1549, 143, 1475, 1077, 1553, 894, 798, 1349, 1885, 1162, 1911, 120, 1110, 1718, 635, 942, 230, 1152, 154, 1215, 1430, 1521, 780, 1833, 1161, 47, 977, 714, 306),		
		--(62, 119, 242, 38, 67, 246, 55, 252, 233, 46, 101, 25, 165, 21, 141, 246, 126, 85, 8, 35, 78, 148, 28, 178, 247, 154, 230, 5, 96, 196, 242, 175, 234, 12, 212, 114, 56, 73, 40, 60, 2, 24, 187, 123, 176, 233, 143, 13, 142, 45, 179, 82, 177, 243, 120, 104, 252, 229, 91, 114, 148, 249, 129, 59, 162, 9, 127, 49, 96, 197, 181, 203, 118, 11, 16, 164, 65, 1, 89, 110, 112, 125, 12, 101, 32, 117, 76, 122, 231, 100, 146, 235, 84, 167, 78, 140, 166, 137, 214, 253, 3, 240, 105, 246, 102, 55, 252, 24, 51, 246, 25, 113, 140, 130, 107, 208, 246, 70, 147, 222, 52, 12, 214, 217, 170, 1, 175, 210, 226, 161, 178, 143, 51, 240, 226, 16, 213, 91, 237, 232, 84, 8, 20, 219, 247, 78, 241, 218, 216, 208, 211, 121, 167, 39, 165, 253, 151, 119, 131, 170, 166, 222, 56, 204, 200, 138, 184, 23, 72, 91, 0, 132, 42, 117, 211, 155, 71, 240, 33, 117, 146, 178, 169, 253, 119, 121, 125, 224, 29, 70, 159, 81, 136, 29, 169, 145, 24, 87, 161, 60, 119, 127, 155, 250, 237, 128, 213, 144, 54, 126, 65, 151, 251, 47, 221, 77, 237, 19, 134, 44, 228, 150, 176, 181, 133, 50, 242, 159, 119, 106, 159, 81, 21, 43, 247, 247, 137, 41, 72, 246, 150, 139, 124, 16, 165, 97, 176, 62, 65, 217, 194, 84, 158, 255, 185, 113, 241, 29, 248, 33, 55, 53, 245, 160, 170, 178, 187, 40, 125, 54, 206, 34, 94, 101, 108, 93, 136, 97, 100, 79, 220, 90, 255, 232, 254, 29, 159, 58, 25, 4, 202, 166, 237, 246, 147, 229, 210, 84, 126, 175, 136, 42, 224, 154, 225, 32, 52, 198, 126, 69, 221, 142, 167, 226, 15, 184, 209, 185, 95, 20, 115, 22, 65, 140, 173, 89, 42, 31, 42, 67, 107, 182, 217, 211, 90, 5, 19, 15, 192, 165, 246, 90, 155, 5, 212, 157, 103, 36, 232, 202, 145, 185, 141, 177, 247, 30, 226, 80, 57, 63, 9, 116, 27, 113, 251, 33, 171, 201, 103, 84, 80, 144, 117, 104, 138, 6, 188, 226, 156, 201, 43, 130, 109, 135, 139, 225, 169, 7, 160, 242, 6, 185, 129, 114, 37, 205, 131, 6, 89, 42, 92, 100, 221, 150, 81, 225, 66, 201, 23, 245, 43, 69, 46, 89, 248, 35, 38, 171, 63, 12, 173, 135, 128, 30, 41, 107, 92, 231, 183, 11, 254, 9, 80, 69, 120, 92, 165, 152, 4, 158, 54, 233, 56, 64, 86, 165, 160, 93, 178, 154, 83, 101, 53, 37, 66, 240, 195, 235, 132, 183, 139, 121, 181, 213, 63, 88, 93, 42, 234, 136, 198, 132, 136, 175, 211, 241, 252, 36, 143, 143, 209, 132, 178, 215, 166, 177, 80, 197, 176, 25, 225, 231, 179, 249, 168, 155, 93, 250, 34, 156, 219, 255, 163, 24, 128, 234, 206, 232, 232, 8, 146, 242, 123, 176, 48, 24, 169, 171, 238, 197, 211, 34, 39, 177, 126, 154, 142, 170, 70, 176, 237, 15, 250, 67, 240, 17, 187, 15, 184, 177, 7, 111, 111, 186, 217, 101, 243, 131, 121, 152, 162, 156, 59, 98, 237, 251, 25, 146, 54, 47, 43, 237, 44, 15, 14, 73, 253, 39, 201, 210, 36, 19, 183, 32, 33, 3, 141, 105, 233, 174, 33, 168, 159, 235, 132, 3, 63, 242, 193, 126, 208, 4, 241, 85, 210, 72, 230, 95, 60, 224, 109, 237, 88, 115, 135, 59, 78, 90, 226, 146, 181, 0, 45, 78, 45, 123, 15, 137),
		(165, 57, 101, 115, 149, 111, 165, 88, 187, 42, 121, 5, 218, 100, 241, 200, 201, 181, 226, 249, 149, 68, 118, 182, 40, 120, 36, 110, 62, 12, 63, 142, 109, 194, 25, 28, 94, 1, 90, 167, 117, 40, 88, 53, 116, 155, 78, 120, 136, 183, 103, 68, 141, 192, 18, 11, 187, 167, 147, 58, 80, 248, 125, 236, 176, 163, 238, 95, 30, 3, 82, 248, 21, 203, 144, 240, 167, 197, 63, 182, 209, 50, 162, 3, 241, 113, 193, 196, 198, 217, 32, 20, 224, 2, 90, 236, 254, 231, 19, 105, 84, 94, 226, 210, 251, 56, 124, 193, 225, 220, 160, 249, 13, 159, 154, 119, 84, 101, 212, 107, 22, 236, 210, 101, 43, 167, 89, 246, 185, 132, 29, 13, 99, 203, 93, 158, 122, 220, 4, 251, 138, 104, 229, 131, 32, 212, 26, 250, 189, 193, 194, 138, 246, 13, 6, 35, 128, 55, 94, 22, 171, 209, 133, 58, 208, 72, 114, 84, 238, 43, 207, 156, 154, 87, 34, 29, 165, 39, 128, 103, 143, 101, 194, 13, 64, 192, 213, 94, 149, 253, 99, 79, 8, 29, 150, 247, 135, 205, 121, 244, 99, 63, 36, 118, 2, 133, 217, 69, 72, 122, 59, 99, 39, 241, 136, 214, 108, 138, 179, 238, 185, 195, 142, 2, 165, 128, 165, 202, 227, 251, 136, 184, 98, 206, 228, 157, 69, 59, 178, 147, 195, 72, 147, 9, 207, 85, 218, 104, 221, 19, 172, 90, 218, 192, 71, 199, 135, 206, 209, 92, 141, 150, 182, 225, 161, 7, 154, 92, 173, 3, 37, 143, 75, 150, 145, 90, 219, 58, 192, 92, 175, 159, 227, 9, 233, 155, 243, 207, 151, 197, 72, 78, 125, 143, 255, 71, 252, 197, 36, 198, 209, 34, 129, 228, 72, 206, 19, 95, 115, 15, 20, 0, 85, 104, 10, 61, 53, 62, 63, 60, 122, 243, 122, 144, 47, 139, 80, 251, 72, 96, 33, 13, 116, 172, 70, 81, 113, 243, 118, 243, 7, 193, 186, 56, 124, 237, 12, 206, 6, 159, 13, 58, 240, 227, 91, 191, 201, 254, 75, 192, 135, 244, 147, 101, 250, 134, 153, 75, 236, 95, 113, 27, 133, 81, 222, 108, 7, 196, 190, 23, 163, 182, 185, 30, 102, 228, 170, 36, 28, 90, 161, 30, 4, 222, 215, 181, 30, 225, 57, 118, 93, 212, 47, 180, 7, 156, 98, 81, 222, 247, 218, 55, 90, 67, 34, 188, 224, 56, 234, 68, 158, 39, 242, 239, 8, 124, 248, 59, 190, 55, 147, 26, 244, 4, 141, 202, 139, 144, 169, 243, 101, 102, 95, 170, 201, 105, 17, 50, 176, 142, 61, 175, 83, 2, 111, 165, 93, 76, 29, 123, 136, 15, 187, 243, 55, 71, 238, 28, 46, 13, 91, 61, 162, 34, 119, 59, 238, 205, 244, 92, 159, 196, 117, 180, 32, 177, 122, 19, 24, 228, 137, 128, 173, 173, 20, 0, 250, 39, 214, 146, 64, 76, 43, 48, 85, 207, 37, 119, 55, 208, 171, 82, 5, 231, 50, 240, 129, 246, 208, 152, 96, 12, 96, 180, 61, 248, 194, 62, 231, 147, 40, 247, 201, 252, 46, 73, 115, 106, 121, 232, 77, 22, 8, 115, 61, 229, 216, 253, 246, 123, 170, 24, 252, 168, 107, 201, 188, 25, 246, 78, 218, 218, 206, 0, 174, 115, 139, 239, 85, 198, 136, 1, 65, 191, 59, 68, 188, 58, 95, 247, 226, 162, 169, 116, 172, 100, 102, 142, 166, 90, 33, 48, 208, 1, 236, 64, 162, 131, 75, 137, 147, 214, 110, 147, 149, 101, 71, 249, 137, 135, 108, 113, 74, 195, 50, 105, 240, 227, 674),
		(0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, 1, 1, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, -1, 0, 0, -1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0),
		"00111100110011001110010111100001101100100001011001101001110110101100101001011111010000111000101111011000011101011111111010000100"
		);
		
        
        --check_dec(
        --(157, 246, 66, 249, 58, 70, 105, 32, 192, 30, 219, 90, 44, 92, 44, 15, 150, 172, 45, 62, 169, 214, 38, 94, 222, 182, 79, 255, 57, 141, 5, 117, 191, 22, 77, 190, 123, 129, 233, 175, 129, 252, 35, 41, 144, 152, 35, 197, 234, 225, 94, 155, 235, 38, 188, 3, 173, 0, 9, 90, 233, 197, 36, 210, 121, 163, 18, 193, 247, 149, 67, 250, 86, 127, 74, 140, 243, 229, 31, 76, 136, 22, 159, 104, 95, 228, 118, 6, 116, 231, 222, 232, 32, 252, 238, 152, 80, 70, 168, 217, 229, 171, 58, 166, 59, 221, 152, 67, 163, 121, 225, 142, 0, 185, 105, 232, 15, 152, 239, 249, 15, 76, 117, 91, 235, 214, 31, 78, 73, 67, 158, 135, 29, 140, 251, 229, 66, 28, 199, 212, 65, 3, 42, 146, 147, 236, 45, 185, 197, 59, 4, 242, 241, 115, 52, 37, 49, 45, 172, 54, 220, 74, 58, 150, 31, 253, 24, 169, 109, 124, 196, 219, 68, 247, 119, 66, 248, 13, 35, 237, 73, 3, 183, 237, 97, 122, 236, 250, 182, 36, 18, 253, 3, 225, 151, 74, 214, 228, 1, 96, 202, 141, 113, 156, 34, 155, 235, 187, 67, 112, 213, 157, 226, 80, 186, 104, 72, 81, 19, 3, 70, 80, 206, 206, 149, 189, 29, 87, 224, 96, 14, 72, 112, 17, 183, 240, 132, 164, 55, 9, 160, 63, 51, 52, 217, 167, 247, 49, 135, 88, 145, 232, 180, 140, 201, 213, 28, 54, 96, 254, 245, 226, 227, 182, 248, 238, 54, 241, 163, 239, 189, 75, 242, 11, 24, 66, 31, 153, 214, 85, 20, 145, 123, 211, 92, 19, 22, 70, 253, 107, 46, 44, 216, 158, 74, 67, 240, 45, 218, 36, 167, 199, 195, 155, 139, 237, 105, 20, 231, 199, 109, 183, 196, 214, 130, 162, 121, 222, 250, 170, 137, 143, 19, 151, 175, 76, 26, 129, 29, 119, 250, 183, 136, 106, 161, 80, 99, 153, 5, 250, 167, 140, 187, 167, 115, 74, 249, 182, 70, 173, 125, 153, 3, 133, 125, 80, 243, 254, 202, 117, 27, 165, 90, 13, 11, 44, 250, 64, 1, 135, 24, 78, 113, 204, 235, 203, 142, 179, 109, 2, 143, 228, 9, 218, 186, 247, 196, 199, 232, 22, 89, 96, 19, 151, 126, 77, 40, 108, 143, 33, 130, 64, 69, 120, 251, 50, 167, 172, 213, 30, 156, 104, 43, 252, 128, 126, 233, 204, 14, 102, 117, 63, 6, 81, 18, 28, 152, 97, 35, 241, 40, 155, 83, 162, 37, 243, 80, 46, 90, 51, 165, 99, 198, 37, 112, 221, 83, 26, 6, 120, 2, 114, 246, 240, 71, 118, 22, 194, 112, 118, 161, 104, 5, 242, 36, 5, 181, 255, 175, 14, 37, 81, 70, 125, 196, 219, 103, 194, 180, 50, 184, 212, 79, 16, 107, 49, 26, 74, 35, 215, 178, 14, 65, 0, 29, 239, 116, 37, 74, 55, 90, 192, 37, 254, 72, 30, 167, 178, 249, 85, 108, 35, 18, 78, 127, 92, 114, 216, 36, 49, 69, 238, 76, 162, 102, 135, 36, 178, 233, 108, 171, 248, 175, 158, 129, 205, 144, 43, 167, 205, 205, 63, 148, 190, 107, 214, 187, 96, 244, 97, 66, 237, 170, 200, 129, 90, 91, 222, 204, 128, 223, 145, 83, 202, 214, 105, 156, 227, 178, 107, 76, 40, 195, 53, 119, 36, 76, 230, 133, 162, 241, 243, 30, 143, 220, 32, 173, 170, 108, 188, 10, 127, 121, 100, 2, 147, 187, 103, 155, 149, 219, 144, 233, 101, 31, 199, 235, 180, 241, 190, 231, 68, 87, 241, 252, 237, 220, 199),
        
        --);
		
		
end process;


--			GG: for i in PolyDegree-1 downto 0 generate
--				PolyA_tmp(i) <= std_logic_vector(to_unsigned(c1(i), LongModLen-1));
--				PolyB_tmp(i) <= std_logic_vector(to_unsigned(c2(i), ShortModLen-1));
--				PolyR_tmp(i) <= std_logic_vector(to_signed(c3(i), 2));
--				
--			end generate GG;




end a1;
