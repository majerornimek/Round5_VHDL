library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
use ieee.numeric_std.all;
use IEEE.math_real.all;


package XEf_constants is  -- R5ND_1KEM_0C

type RTab is array(natural range<>) of std_logic_vector(63 downto 0);
type BitTab is array(natural range<>) of std_logic_vector(7 downto 0);

type wt is array(0 to 255, 0 to 10) of integer;

constant wire_tab : wt :=
(
(0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0),
(0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1),
(0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2),
(0, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3),
(0, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4),
(0, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5),
(0, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6),
(0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7),
(0, 8, 8, 8, 8, 8, 8, 8, 8, 8, 0),
(0, 9, 9, 9, 9, 9, 9, 9, 9, 9, 1),
(0, 10, 10, 10, 10, 10, 10, 10, 10, 10, 2),
(0, 11, 11, 11, 11, 11, 11, 11, 11, 11, 3),
(0, 12, 12, 12, 12, 12, 12, 12, 12, 12, 4),
(0, 13, 13, 13, 13, 13, 13, 13, 13, 13, 5),
(0, 14, 14, 14, 14, 14, 14, 14, 14, 14, 6),
(0, 15, 15, 15, 15, 15, 15, 15, 15, 15, 7),
(1, 0, 16, 16, 16, 16, 16, 16, 16, 16, 0),
(1, 1, 0, 17, 17, 17, 17, 17, 17, 17, 1),
(1, 2, 1, 18, 18, 18, 18, 18, 18, 18, 2),
(1, 3, 2, 0, 19, 19, 19, 19, 19, 19, 3),
(1, 4, 3, 1, 20, 20, 20, 20, 20, 20, 4),
(1, 5, 4, 2, 0, 21, 21, 21, 21, 21, 5),
(1, 6, 5, 3, 1, 22, 22, 22, 22, 22, 6),
(1, 7, 6, 4, 2, 0, 23, 23, 23, 23, 7),
(1, 8, 7, 5, 3, 1, 24, 24, 24, 24, 0),
(1, 9, 8, 6, 4, 2, 0, 25, 25, 25, 1),
(1, 10, 9, 7, 5, 3, 1, 26, 26, 26, 2),
(1, 11, 10, 8, 6, 4, 2, 27, 27, 27, 3),
(1, 12, 11, 9, 7, 5, 3, 28, 28, 28, 4),
(1, 13, 12, 10, 8, 6, 4, 0, 29, 29, 5),
(1, 14, 13, 11, 9, 7, 5, 1, 30, 30, 6),
(1, 15, 14, 12, 10, 8, 6, 2, 0, 31, 7),
(2, 0, 15, 13, 11, 9, 7, 3, 1, 32, 0),
(2, 1, 16, 14, 12, 10, 8, 4, 2, 33, 1),
(2, 2, 0, 15, 13, 11, 9, 5, 3, 34, 2),
(2, 3, 1, 16, 14, 12, 10, 6, 4, 35, 3),
(2, 4, 2, 17, 15, 13, 11, 7, 5, 36, 4),
(2, 5, 3, 18, 16, 14, 12, 8, 6, 0, 5),
(2, 6, 4, 0, 17, 15, 13, 9, 7, 1, 6),
(2, 7, 5, 1, 18, 16, 14, 10, 8, 2, 7),
(2, 8, 6, 2, 19, 17, 15, 11, 9, 3, 0),
(2, 9, 7, 3, 20, 18, 16, 12, 10, 4, 1),
(2, 10, 8, 4, 0, 19, 17, 13, 11, 5, 2),
(2, 11, 9, 5, 1, 20, 18, 14, 12, 6, 3),
(2, 12, 10, 6, 2, 21, 19, 15, 13, 7, 4),
(2, 13, 11, 7, 3, 22, 20, 16, 14, 8, 5),
(2, 14, 12, 8, 4, 0, 21, 17, 15, 9, 6),
(2, 15, 13, 9, 5, 1, 22, 18, 16, 10, 7),
(3, 0, 14, 10, 6, 2, 23, 19, 17, 11, 0),
(3, 1, 15, 11, 7, 3, 24, 20, 18, 12, 1),
(3, 2, 16, 12, 8, 4, 0, 21, 19, 13, 2),
(3, 3, 0, 13, 9, 5, 1, 22, 20, 14, 3),
(3, 4, 1, 14, 10, 6, 2, 23, 21, 15, 4),
(3, 5, 2, 15, 11, 7, 3, 24, 22, 16, 5),
(3, 6, 3, 16, 12, 8, 4, 25, 23, 17, 6),
(3, 7, 4, 17, 13, 9, 5, 26, 24, 18, 7),
(3, 8, 5, 18, 14, 10, 6, 27, 25, 19, 0),
(3, 9, 6, 0, 15, 11, 7, 28, 26, 20, 1),
(3, 10, 7, 1, 16, 12, 8, 0, 27, 21, 2),
(3, 11, 8, 2, 17, 13, 9, 1, 28, 22, 3),
(3, 12, 9, 3, 18, 14, 10, 2, 29, 23, 4),
(3, 13, 10, 4, 19, 15, 11, 3, 30, 24, 5),
(3, 14, 11, 5, 20, 16, 12, 4, 0, 25, 6),
(3, 15, 12, 6, 0, 17, 13, 5, 1, 26, 7),
(4, 0, 13, 7, 1, 18, 14, 6, 2, 27, 0),
(4, 1, 14, 8, 2, 19, 15, 7, 3, 28, 1),
(4, 2, 15, 9, 3, 20, 16, 8, 4, 29, 2),
(4, 3, 16, 10, 4, 21, 17, 9, 5, 30, 3),
(4, 4, 0, 11, 5, 22, 18, 10, 6, 31, 4),
(4, 5, 1, 12, 6, 0, 19, 11, 7, 32, 5),
(4, 6, 2, 13, 7, 1, 20, 12, 8, 33, 6),
(4, 7, 3, 14, 8, 2, 21, 13, 9, 34, 7),
(4, 8, 4, 15, 9, 3, 22, 14, 10, 35, 0),
(4, 9, 5, 16, 10, 4, 23, 15, 11, 36, 1),
(4, 10, 6, 17, 11, 5, 24, 16, 12, 0, 2),
(4, 11, 7, 18, 12, 6, 0, 17, 13, 1, 3),
(4, 12, 8, 0, 13, 7, 1, 18, 14, 2, 4),
(4, 13, 9, 1, 14, 8, 2, 19, 15, 3, 5),
(4, 14, 10, 2, 15, 9, 3, 20, 16, 4, 6),
(4, 15, 11, 3, 16, 10, 4, 21, 17, 5, 7),
(5, 0, 12, 4, 17, 11, 5, 22, 18, 6, 0),
(5, 1, 13, 5, 18, 12, 6, 23, 19, 7, 1),
(5, 2, 14, 6, 19, 13, 7, 24, 20, 8, 2),
(5, 3, 15, 7, 20, 14, 8, 25, 21, 9, 3),
(5, 4, 16, 8, 0, 15, 9, 26, 22, 10, 4),
(5, 5, 0, 9, 1, 16, 10, 27, 23, 11, 5),
(5, 6, 1, 10, 2, 17, 11, 28, 24, 12, 6),
(5, 7, 2, 11, 3, 18, 12, 0, 25, 13, 7),
(5, 8, 3, 12, 4, 19, 13, 1, 26, 14, 0),
(5, 9, 4, 13, 5, 20, 14, 2, 27, 15, 1),
(5, 10, 5, 14, 6, 21, 15, 3, 28, 16, 2),
(5, 11, 6, 15, 7, 22, 16, 4, 29, 17, 3),
(5, 12, 7, 16, 8, 0, 17, 5, 30, 18, 4),
(5, 13, 8, 17, 9, 1, 18, 6, 0, 19, 5),
(5, 14, 9, 18, 10, 2, 19, 7, 1, 20, 6),
(5, 15, 10, 0, 11, 3, 20, 8, 2, 21, 7),
(6, 0, 11, 1, 12, 4, 21, 9, 3, 22, 0),
(6, 1, 12, 2, 13, 5, 22, 10, 4, 23, 1),
(6, 2, 13, 3, 14, 6, 23, 11, 5, 24, 2),
(6, 3, 14, 4, 15, 7, 24, 12, 6, 25, 3),
(6, 4, 15, 5, 16, 8, 0, 13, 7, 26, 4),
(6, 5, 16, 6, 17, 9, 1, 14, 8, 27, 5),
(6, 6, 0, 7, 18, 10, 2, 15, 9, 28, 6),
(6, 7, 1, 8, 19, 11, 3, 16, 10, 29, 7),
(6, 8, 2, 9, 20, 12, 4, 17, 11, 30, 0),
(6, 9, 3, 10, 0, 13, 5, 18, 12, 31, 1),
(6, 10, 4, 11, 1, 14, 6, 19, 13, 32, 2),
(6, 11, 5, 12, 2, 15, 7, 20, 14, 33, 3),
(6, 12, 6, 13, 3, 16, 8, 21, 15, 34, 4),
(6, 13, 7, 14, 4, 17, 9, 22, 16, 35, 5),
(6, 14, 8, 15, 5, 18, 10, 23, 17, 36, 6),
(6, 15, 9, 16, 6, 19, 11, 24, 18, 0, 7),
(7, 0, 10, 17, 7, 20, 12, 25, 19, 1, 0),
(7, 1, 11, 18, 8, 21, 13, 26, 20, 2, 1),
(7, 2, 12, 0, 9, 22, 14, 27, 21, 3, 2),
(7, 3, 13, 1, 10, 0, 15, 28, 22, 4, 3),
(7, 4, 14, 2, 11, 1, 16, 0, 23, 5, 4),
(7, 5, 15, 3, 12, 2, 17, 1, 24, 6, 5),
(7, 6, 16, 4, 13, 3, 18, 2, 25, 7, 6),
(7, 7, 0, 5, 14, 4, 19, 3, 26, 8, 7),
(7, 8, 1, 6, 15, 5, 20, 4, 27, 9, 0),
(7, 9, 2, 7, 16, 6, 21, 5, 28, 10, 1),
(7, 10, 3, 8, 17, 7, 22, 6, 29, 11, 2),
(7, 11, 4, 9, 18, 8, 23, 7, 30, 12, 3),
(7, 12, 5, 10, 19, 9, 24, 8, 0, 13, 4),
(7, 13, 6, 11, 20, 10, 0, 9, 1, 14, 5),
(7, 14, 7, 12, 0, 11, 1, 10, 2, 15, 6),
(7, 15, 8, 13, 1, 12, 2, 11, 3, 16, 7),
(8, 0, 9, 14, 2, 13, 3, 12, 4, 17, 0),
(8, 1, 10, 15, 3, 14, 4, 13, 5, 18, 1),
(8, 2, 11, 16, 4, 15, 5, 14, 6, 19, 2),
(8, 3, 12, 17, 5, 16, 6, 15, 7, 20, 3),
(8, 4, 13, 18, 6, 17, 7, 16, 8, 21, 4),
(8, 5, 14, 0, 7, 18, 8, 17, 9, 22, 5),
(8, 6, 15, 1, 8, 19, 9, 18, 10, 23, 6),
(8, 7, 16, 2, 9, 20, 10, 19, 11, 24, 7),
(8, 8, 0, 3, 10, 21, 11, 20, 12, 25, 0),
(8, 9, 1, 4, 11, 22, 12, 21, 13, 26, 1),
(8, 10, 2, 5, 12, 0, 13, 22, 14, 27, 2),
(8, 11, 3, 6, 13, 1, 14, 23, 15, 28, 3),
(8, 12, 4, 7, 14, 2, 15, 24, 16, 29, 4),
(8, 13, 5, 8, 15, 3, 16, 25, 17, 30, 5),
(8, 14, 6, 9, 16, 4, 17, 26, 18, 31, 6),
(8, 15, 7, 10, 17, 5, 18, 27, 19, 32, 7),
(9, 0, 8, 11, 18, 6, 19, 28, 20, 33, 0),
(9, 1, 9, 12, 19, 7, 20, 0, 21, 34, 1),
(9, 2, 10, 13, 20, 8, 21, 1, 22, 35, 2),
(9, 3, 11, 14, 0, 9, 22, 2, 23, 36, 3),
(9, 4, 12, 15, 1, 10, 23, 3, 24, 0, 4),
(9, 5, 13, 16, 2, 11, 24, 4, 25, 1, 5),
(9, 6, 14, 17, 3, 12, 0, 5, 26, 2, 6),
(9, 7, 15, 18, 4, 13, 1, 6, 27, 3, 7),
(9, 8, 16, 0, 5, 14, 2, 7, 28, 4, 0),
(9, 9, 0, 1, 6, 15, 3, 8, 29, 5, 1),
(9, 10, 1, 2, 7, 16, 4, 9, 30, 6, 2),
(9, 11, 2, 3, 8, 17, 5, 10, 0, 7, 3),
(9, 12, 3, 4, 9, 18, 6, 11, 1, 8, 4),
(9, 13, 4, 5, 10, 19, 7, 12, 2, 9, 5),
(9, 14, 5, 6, 11, 20, 8, 13, 3, 10, 6),
(9, 15, 6, 7, 12, 21, 9, 14, 4, 11, 7),
(10, 0, 7, 8, 13, 22, 10, 15, 5, 12, 0),
(10, 1, 8, 9, 14, 0, 11, 16, 6, 13, 1),
(10, 2, 9, 10, 15, 1, 12, 17, 7, 14, 2),
(10, 3, 10, 11, 16, 2, 13, 18, 8, 15, 3),
(10, 4, 11, 12, 17, 3, 14, 19, 9, 16, 4),
(10, 5, 12, 13, 18, 4, 15, 20, 10, 17, 5),
(10, 6, 13, 14, 19, 5, 16, 21, 11, 18, 6),
(10, 7, 14, 15, 20, 6, 17, 22, 12, 19, 7),
(10, 8, 15, 16, 0, 7, 18, 23, 13, 20, 0),
(10, 9, 16, 17, 1, 8, 19, 24, 14, 21, 1),
(10, 10, 0, 18, 2, 9, 20, 25, 15, 22, 2),
(10, 11, 1, 0, 3, 10, 21, 26, 16, 23, 3),
(10, 12, 2, 1, 4, 11, 22, 27, 17, 24, 4),
(10, 13, 3, 2, 5, 12, 23, 28, 18, 25, 5),
(10, 14, 4, 3, 6, 13, 24, 0, 19, 26, 6),
(10, 15, 5, 4, 7, 14, 0, 1, 20, 27, 7),
(11, 0, 6, 5, 8, 15, 1, 2, 21, 28, 0),
(11, 1, 7, 6, 9, 16, 2, 3, 22, 29, 1),
(11, 2, 8, 7, 10, 17, 3, 4, 23, 30, 2),
(11, 3, 9, 8, 11, 18, 4, 5, 24, 31, 3),
(11, 4, 10, 9, 12, 19, 5, 6, 25, 32, 4),
(11, 5, 11, 10, 13, 20, 6, 7, 26, 33, 5),
(11, 6, 12, 11, 14, 21, 7, 8, 27, 34, 6),
(11, 7, 13, 12, 15, 22, 8, 9, 28, 35, 7),
(11, 8, 14, 13, 16, 0, 9, 10, 29, 36, 0),
(11, 9, 15, 14, 17, 1, 10, 11, 30, 0, 1),
(11, 10, 16, 15, 18, 2, 11, 12, 0, 1, 2),
(11, 11, 0, 16, 19, 3, 12, 13, 1, 2, 3),
(11, 12, 1, 17, 20, 4, 13, 14, 2, 3, 4),
(11, 13, 2, 18, 0, 5, 14, 15, 3, 4, 5),
(11, 14, 3, 0, 1, 6, 15, 16, 4, 5, 6),
(11, 15, 4, 1, 2, 7, 16, 17, 5, 6, 7),
(12, 0, 5, 2, 3, 8, 17, 18, 6, 7, 0),
(12, 1, 6, 3, 4, 9, 18, 19, 7, 8, 1),
(12, 2, 7, 4, 5, 10, 19, 20, 8, 9, 2),
(12, 3, 8, 5, 6, 11, 20, 21, 9, 10, 3),
(12, 4, 9, 6, 7, 12, 21, 22, 10, 11, 4),
(12, 5, 10, 7, 8, 13, 22, 23, 11, 12, 5),
(12, 6, 11, 8, 9, 14, 23, 24, 12, 13, 6),
(12, 7, 12, 9, 10, 15, 24, 25, 13, 14, 7),
(12, 8, 13, 10, 11, 16, 0, 26, 14, 15, 0),
(12, 9, 14, 11, 12, 17, 1, 27, 15, 16, 1),
(12, 10, 15, 12, 13, 18, 2, 28, 16, 17, 2),
(12, 11, 16, 13, 14, 19, 3, 0, 17, 18, 3),
(12, 12, 0, 14, 15, 20, 4, 1, 18, 19, 4),
(12, 13, 1, 15, 16, 21, 5, 2, 19, 20, 5),
(12, 14, 2, 16, 17, 22, 6, 3, 20, 21, 6),
(12, 15, 3, 17, 18, 0, 7, 4, 21, 22, 7),
(13, 0, 4, 18, 19, 1, 8, 5, 22, 23, 0),
(13, 1, 5, 0, 20, 2, 9, 6, 23, 24, 1),
(13, 2, 6, 1, 0, 3, 10, 7, 24, 25, 2),
(13, 3, 7, 2, 1, 4, 11, 8, 25, 26, 3),
(13, 4, 8, 3, 2, 5, 12, 9, 26, 27, 4),
(13, 5, 9, 4, 3, 6, 13, 10, 27, 28, 5),
(13, 6, 10, 5, 4, 7, 14, 11, 28, 29, 6),
(13, 7, 11, 6, 5, 8, 15, 12, 29, 30, 7),
(13, 8, 12, 7, 6, 9, 16, 13, 30, 31, 0),
(13, 9, 13, 8, 7, 10, 17, 14, 0, 32, 1),
(13, 10, 14, 9, 8, 11, 18, 15, 1, 33, 2),
(13, 11, 15, 10, 9, 12, 19, 16, 2, 34, 3),
(13, 12, 16, 11, 10, 13, 20, 17, 3, 35, 4),
(13, 13, 0, 12, 11, 14, 21, 18, 4, 36, 5),
(13, 14, 1, 13, 12, 15, 22, 19, 5, 0, 6),
(13, 15, 2, 14, 13, 16, 23, 20, 6, 1, 7),
(14, 0, 3, 15, 14, 17, 24, 21, 7, 2, 0),
(14, 1, 4, 16, 15, 18, 0, 22, 8, 3, 1),
(14, 2, 5, 17, 16, 19, 1, 23, 9, 4, 2),
(14, 3, 6, 18, 17, 20, 2, 24, 10, 5, 3),
(14, 4, 7, 0, 18, 21, 3, 25, 11, 6, 4),
(14, 5, 8, 1, 19, 22, 4, 26, 12, 7, 5),
(14, 6, 9, 2, 20, 0, 5, 27, 13, 8, 6),
(14, 7, 10, 3, 0, 1, 6, 28, 14, 9, 7),
(14, 8, 11, 4, 1, 2, 7, 0, 15, 10, 0),
(14, 9, 12, 5, 2, 3, 8, 1, 16, 11, 1),
(14, 10, 13, 6, 3, 4, 9, 2, 17, 12, 2),
(14, 11, 14, 7, 4, 5, 10, 3, 18, 13, 3),
(14, 12, 15, 8, 5, 6, 11, 4, 19, 14, 4),
(14, 13, 16, 9, 6, 7, 12, 5, 20, 15, 5),
(14, 14, 0, 10, 7, 8, 13, 6, 21, 16, 6),
(14, 15, 1, 11, 8, 9, 14, 7, 22, 17, 7),
(15, 0, 2, 12, 9, 10, 15, 8, 23, 18, 0),
(15, 1, 3, 13, 10, 11, 16, 9, 24, 19, 1),
(15, 2, 4, 14, 11, 12, 17, 10, 25, 20, 2),
(15, 3, 5, 15, 12, 13, 18, 11, 26, 21, 3),
(15, 4, 6, 16, 13, 14, 19, 12, 27, 22, 4),
(15, 5, 7, 17, 14, 15, 20, 13, 28, 23, 5),
(15, 6, 8, 18, 15, 16, 21, 14, 29, 24, 6),
(15, 7, 9, 0, 16, 17, 22, 15, 30, 25, 7),
(15, 8, 10, 1, 17, 18, 23, 16, 0, 26, 0),
(15, 9, 11, 2, 18, 19, 24, 17, 1, 27, 1),
(15, 10, 12, 3, 19, 20, 0, 18, 2, 28, 2),
(15, 11, 13, 4, 20, 21, 1, 19, 3, 29, 3),
(15, 12, 14, 5, 0, 22, 2, 20, 4, 30, 4),
(15, 13, 15, 6, 1, 0, 3, 21, 5, 31, 5),
(15, 14, 16, 7, 2, 1, 4, 22, 6, 32, 6),
(15, 15, 0, 8, 3, 2, 5, 23, 7, 33, 7)
-- (std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(25,6)), std_logic_vector(to_unsigned(25,6)), std_logic_vector(to_unsigned(25,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(26,6)), std_logic_vector(to_unsigned(26,6)), std_logic_vector(to_unsigned(26,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(27,6)), std_logic_vector(to_unsigned(27,6)), std_logic_vector(to_unsigned(27,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(28,6)), std_logic_vector(to_unsigned(28,6)), std_logic_vector(to_unsigned(28,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(29,6)), std_logic_vector(to_unsigned(29,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(30,6)), std_logic_vector(to_unsigned(30,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(31,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(32,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(33,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(34,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(35,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(36,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(25,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(26,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(27,6)), std_logic_vector(to_unsigned(25,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(28,6)), std_logic_vector(to_unsigned(26,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(27,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(28,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(29,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(30,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(25,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(26,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(27,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(28,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(29,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(30,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(31,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(32,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(33,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(34,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(35,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(36,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(25,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(26,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(27,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(28,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(25,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(26,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(27,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(28,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(29,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(30,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(25,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(26,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(27,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(28,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(29,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(30,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(31,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(32,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(33,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(34,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(35,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(36,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(25,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(26,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(27,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(28,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(25,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(26,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(27,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(28,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(29,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(30,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(25,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(26,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(27,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(28,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(29,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(25,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(30,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(26,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(31,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(27,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(32,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(28,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(33,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(34,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(35,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(36,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(25,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(26,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(27,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(28,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(29,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(30,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(25,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(26,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(27,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(28,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(25,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(26,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(27,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(28,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(29,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(30,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(31,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(25,6)), std_logic_vector(to_unsigned(32,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(26,6)), std_logic_vector(to_unsigned(33,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(27,6)), std_logic_vector(to_unsigned(34,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(28,6)), std_logic_vector(to_unsigned(35,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(29,6)), std_logic_vector(to_unsigned(36,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(30,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(25,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(26,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(27,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(28,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(25,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(25,6)), std_logic_vector(to_unsigned(26,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(26,6)), std_logic_vector(to_unsigned(27,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(27,6)), std_logic_vector(to_unsigned(28,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(28,6)), std_logic_vector(to_unsigned(29,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(29,6)), std_logic_vector(to_unsigned(30,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(30,6)), std_logic_vector(to_unsigned(31,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(32,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(33,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(34,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(35,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(36,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(25,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(26,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(27,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(28,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(25,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(26,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(27,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(28,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(29,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(30,6)), std_logic_vector(to_unsigned(25,6)), std_logic_vector(to_unsigned(7,6))),
-- (std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(26,6)), std_logic_vector(to_unsigned(0,6))),
-- (std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(9,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(24,6)), std_logic_vector(to_unsigned(17,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(27,6)), std_logic_vector(to_unsigned(1,6))),
-- (std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(10,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(18,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(28,6)), std_logic_vector(to_unsigned(2,6))),
-- (std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(11,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(19,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(29,6)), std_logic_vector(to_unsigned(3,6))),
-- (std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(12,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(20,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(30,6)), std_logic_vector(to_unsigned(4,6))),
-- (std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(13,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(21,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(31,6)), std_logic_vector(to_unsigned(5,6))),
-- (std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(14,6)), std_logic_vector(to_unsigned(16,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(1,6)), std_logic_vector(to_unsigned(4,6)), std_logic_vector(to_unsigned(22,6)), std_logic_vector(to_unsigned(6,6)), std_logic_vector(to_unsigned(32,6)), std_logic_vector(to_unsigned(6,6))),
-- (std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(15,6)), std_logic_vector(to_unsigned(0,6)), std_logic_vector(to_unsigned(8,6)), std_logic_vector(to_unsigned(3,6)), std_logic_vector(to_unsigned(2,6)), std_logic_vector(to_unsigned(5,6)), std_logic_vector(to_unsigned(23,6)), std_logic_vector(to_unsigned(7,6)), std_logic_vector(to_unsigned(33,6)), std_logic_vector(to_unsigned(7,6)))
);

end package;
