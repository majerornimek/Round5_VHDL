library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
use ieee.numeric_std.all;

library work;
use work.Round5_constants.all;

entity Mul_Poly_TB is
end entity; 

architecture a1 of Mul_Poly_TB is 
component Mul_Poly is 
	port (
		PolyA	: in NTRUPoly(PolyDegree downto 0);
		PolyB	: in Trinomial(PolyDegree downto 0); 
		clk		: in std_logic;
		Start	: in std_logic;
		Rst		: in std_logic;
		OpType	: in std_logic;
		Done	: out std_logic;
		LongRes	: out NTRUPoly(PolyDegree downto 0);
		ShortRes: out ShortPoly(PolyDegree downto 0)
	);
end component;
signal inA, outC : NTRUPoly(PolyDegree downto 0);
signal inB : Trinomial(PolyDegree downto  0); 
signal outS : ShortPoly(PolyDegree downto  0);
signal clk, start_tmp, rst_tmp, op_tmp, done_tmp : std_logic;
constant CLK_PERIOD : time := 10 ps;
type input_array is array(PolyDegree downto 0) of integer;

begin

 clk_process :process
   begin
        clk <= '0';
        wait for CLK_PERIOD/2;  --for half of clock period clk stays at '0'.
        clk <= '1';
        wait for CLK_PERIOD/2;  --for next half of clock period clk stays at '1'.
   end process;
   
   uut: Mul_Poly port map(
    	PolyA	=> inA,
		PolyB	=> inB,
		clk		=> clk,
		Start	=> start_tmp,
		Rst		=> rst_tmp,
		OpType	=> op_tmp,
		Done	=> done_tmp,
		LongRes	=> outC,
		ShortRes=> outS
   );
   
process
	
	procedure check_poly_mul( 	constant PolyA	: in input_array; -- v1
								constant PolyB 	: in input_array; -- v2
								constant typ	: in std_logic; -- norm of v1
								constant res_ex	: in input_array) is
		variable res: input_array;
	begin
		GG: for i in PolyDegree downto 0 loop
			inA(i) <= std_logic_vector(to_signed(PolyA(i), LongModLen-1));
			inB(i) <= std_logic_vector(to_signed(PolyB(i), 2));
		end loop GG; 
		
		wait for CLK_PERIOD;
		rst_tmp <= '1';
		op_tmp <= typ;
		wait for CLK_PERIOD;
		rst_tmp <= '0';
		start_tmp <= '1';
		wait for CLK_PERIOD*700;
		start_tmp <= '0';
		wait for CLK_PERIOD;
		
--		RR: for i in NUM_OF_ELEMENTS-1 downto 0 loop
--			res(i) = to_integer(signed(outC(i)));
--		end loop RR;
--		assert res = res_ex
--		report 	"Unexpected result: " --&
----				"IN1 = " & integer'image(in1) & "; " &
----				"IN2 = " & integer'image(in2) & "; " &
----				"MUL = " & integer'image(res) & "; " &
----				"MUL_expected = " & integer'image(res_ex)
--		severity error;
	end procedure check_poly_mul;
	
	
begin
	
    check_poly_mul((784,2028,1705,574,571,1226,1324,236,642,1876,105,1158,388,1119,1563,204,1977,1595,1048,1785,1845,1345,1894,1990,1591,1753,1276,1568,104,1220,651,511,38,1343,701,1517,402,1727,291,438,381,101,506,35,120,1370,806,362,953,1959,805,606,457,13,1037,1904,614,1745,703,2027,813,1634,2017,917,1269,910,717,497,1325,2017,1869,266,992,1904,204,1208,1363,801,799,1535,965,1104,253,1493,1360,122,1850,1903,1775,1021,972,1961,1545,1390,255,595,1105,1037,937,689,802,1039,1930,1728,134,1894,1650,1230,294,1382,651,1966,1544,459,947,1983,491,648,1363,2040,279,50,880,700,301,816,319,934,1204,263,1196,1348,1395,1059,1238,942,69,1105,319,266,1794,1591,1264,439,1462,1244,1812,1404,1920,153,653,61,299,411,1528,404,745,12,894,1573,961,1716,1725,863,1623,906,1992,188,1297,1113,1829,573,949,627,1733,1247,739,777,1926,1765,1630,991,1574,1567,5,1955,693,19,1594,424,509,1947,1761,1201,263,1565,119,1736,1755,349,784,447,1495,455,400,1636,1731,702,1610,1959,964,1396,1673,1970,443,303,1369,959,574,809,719,1659,771,1709,1756,1421,1992,672,1648,792,189,1181,275,466,1171,153,1101,354,969,348,1217,1452,2043,734,1930,1056,1042,1218,218,1313,362,43,945,825,332,1334,707,23,283,904,779,1830,404,1772,1677,1933,574,352,98,762,1384,1433,1717,1455,512,528,1423,435,693,856,116,659,381,129,308,1242,373,86,735,1841,995,1278,1563,669,485,147,1043,2026,1648,1615,934,186,616,2008,1698,314,963,699,148,1271,538,1037,968,947,606,822,1944,1053,1498,1765,1974,1310,352,790,411,1743,1529,142,1514,565,1190,450,164,487,1135,733,15,626,545,1039,828,678,1350,727,791,1909,1314,660,1223,1209,1097,448,1467,603,1352,1836,1854,360,1668,212,1403,1227,461,411,2031,408,1115,38,554,874,1916,1858,2033,1777,1754,1542,1220,1704,1645,1040,366,1279,864,15,932,570,796,692,1342,99,877,713,9,1474,267,501,175,1612,769,1877,831,870,888,1656,231,129,987,560,1611,1828,113,621,1370,786,272,677,718,419,1141,1029,622,549,277,1003,1500,1876,487,320,1429,951,365,1899,138,1162,1625,863,1848,735,15,187,1288,317,1019,663,1591,1987,597,1654,296,1519,1277,1099,954,1891,1904,935,910,2045,149,1735,679,507,1125,221,75,1016,1541,656,750,1717,1585,212,1035,1965,328,1263,1054,1634,968,1512,1269,1334,2045,1783,1306,268,971,1649,126,572,1118,186,1574,1623,1048,1451,289,1785,1563,999,1053,1007,547,586,291,1690,211,255,409,647,325,1951,676,995,59,1841,1239,1026,1509,141,224,772,520,376,125,1039,1598,1141,159,1931,79,1709,1349,475,132,1109,705,916,1261,1331,316,22,904,1670,955,1764,276,285,385,1525,457,823,1392,478,1557,1382,23,1165,500,1272,564,393,442,138,1891,1513,1405,1982,175,895,701,1022,1828,981,50,846,489,1668,885,477,175,991,1089,728,640,724,247,950,1930,644,2016,1174,1857,1061,239,1819,1809,1529,1391,1062,523,1469,1849,154,291,1939,1672,912,1682,840,1730,89,300,1405,1288,374,1021,985,0),
    (0,0,0,0,0,0,0,-1,0,0,0,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,1,0,0,1,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,1,-1,0,0,0,-1,0,0,-1,0,0,0,0,0,0,0,1,0,1,0,0,1,0,0,0,0,0,0,0,-1,1,1,0,0,0,0,0,1,0,0,0,0,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,0,0,0,0,0,0,-1,0,0,0,0,0,0,1,0,0,1,0,0,0,1,0,0,0,0,0,0,0,0,0,0,-1,1,-1,0,0,0,0,0,1,0,0,-1,0,0,0,0,0,0,0,0,0,1,-1,0,1,0,0,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,0,0,0,0,-1,0,-1,0,0,0,1,-1,0,0,0,0,0,0,0,0,-1,0,-1,0,0,0,0,0,-1,0,0,0,0,0,-1,0,0,1,0,0,0,0,0,0,0,0,0,0,-1,0,1,1,0,0,0,0,0,0,0,0,0,0,-1,-1,1,1,0,0,0,0,0,0,1,0,0,-1,-1,0,0,0,0,0,0,1,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,-1,0,0,0,-1,0,0,1,0,0,0,0,1,0,0,0,0,0,0,0,0,0,-1,0,1,0,0,0,0,0,0,0,1,0,0,0,-1,1,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,0,0,1,1,0,0,0,0,0,0,0,-1,0,0,1,1,0,0,0,0,0,0,0,1,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,0,0,0,0,0,0,0,0,0,0,-1,0,0,-1,0,0,-1,0,0,0,0,-1,1,-1,0,0,0,0,0,0,0,-1,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,1,0,0,0,0,0,0,0,0,0,0,-1,0,-1,-1,0,1,0,0,0,0,0,0,0,0,0,0,1,0,1,1,-1,-1,0,0,0,0,0,0,-1,0,0,0,0,0,0,0,0,1,0,0,0,0,-1,0,0,0,0),
   '1',
   (486, 251, 2019, 423, 1295, 1109, 1045, 1240, 366, 353, 1411, 1238, 1126, 1145, 362, 1101, 2022, 1173, 270, 238, 588, 580, 698, 951, 842, 1174, 508, 545, 852, 1539, 1571, 1834, 590, 1536, 1172, 1849, 1059, 918, 1194, 667, 993, 1163, 916, 107, 722, 1319, 1750, 1950, 808, 716, 1849, 1077, 1229, 691, 979, 245, 215, 121, 1943, 1839, 711, 209, 1964, 1533, 1852, 1612, 1021, 1839, 853, 1309, 1540, 1177, 936, 80, 284, 359, 1899, 377, 6, 1214, 794, 899, 1034, 926, 926, 1941, 1163, 1264, 1544, 1163, 1123, 994, 675, 1890, 132, 763, 830, 892, 669, 1608, 502, 1717, 1309, 1385, 394, 696, 763, 1636, 827, 1000, 708, 1437, 1131, 1351, 621, 1801, 1063, 706, 672, 1703, 1848, 2033, 540, 554, 1006, 1725, 1514, 843, 299, 2010, 614, 1143, 1766, 1185, 820, 185, 168, 1023, 579, 1649, 356, 1586, 1804, 84, 969, 518, 113, 1920, 1324, 615, 1976, 299, 189, 1402, 436, 1085, 1088, 1534, 1247, 550, 2012, 857, 1161, 1356, 172, 784, 1650, 522, 377, 433, 1741, 106, 1094, 10, 1685, 1666, 289, 1070, 751, 1715, 390, 771, 590, 807, 1173, 596, 441, 239, 322, 1023, 991, 232, 770, 1529, 229, 283, 962, 70, 1830, 1261, 1515, 1756, 386, 1268, 1528, 458, 383, 1119, 133, 113, 703, 1848, 769, 536, 1588, 1355, 305, 928, 696, 766, 324, 237, 1786, 2025, 1227, 383, 1511, 1504, 1973, 1730, 1845, 991, 920, 966, 211, 844, 1726, 1394, 1618, 1100, 1086, 1782, 1365, 1304, 1029, 1593, 716, 1693, 694, 1143, 1365, 1667, 1801, 673, 1941, 1781, 1050, 525, 355, 1407, 1681, 66, 1997, 1898, 1160, 493, 1503, 808, 978, 356, 993, 81, 6, 1305, 704, 536, 1947, 1970, 445, 1614, 1745, 256, 417, 1190, 693, 1496, 847, 1490, 1529, 134, 997, 1127, 629, 1466, 409, 1786, 173, 1999, 289, 66, 168, 1003, 1688, 47, 1715, 1439, 716, 1231, 1817, 1777, 1905, 736, 681, 188, 1251, 448, 89, 706, 1961, 2014, 604, 1187, 1649, 836, 1223, 336, 172, 858, 2016, 2017, 351, 37, 2027, 1280, 109, 1115, 1043, 1335, 454, 17, 1665, 1501, 1363, 1151, 1522, 2022, 304, 882, 2011, 425, 1136, 73, 90, 1930, 999, 998, 1340, 669, 52, 714, 1922, 1646, 1561, 1142, 145, 1971, 1544, 1571, 842, 1413, 1670, 1641, 1847, 216, 814, 1, 1259, 637, 115, 1542, 2036, 1818, 9, 1311, 1233, 1903, 371, 1686, 1642, 72, 1336, 414, 1626, 1656, 539, 835, 144, 1629, 993, 1117, 1829, 1266, 1094, 379, 2012, 799, 2041, 59, 2027, 1450, 618, 110, 1756, 398, 408, 1783, 873, 1970, 1030, 1177, 1916, 1643, 1079, 1816, 609, 1560, 258, 1303, 1164, 1126, 828, 1108, 164, 908, 995, 1000, 179, 1087, 1682, 1479, 2018, 1015, 561, 1143, 3, 1506, 677, 565, 478, 837, 205, 324, 277, 864, 1368, 348, 1085, 1302, 1516, 136, 445, 547, 655, 271, 423, 778, 1136, 802, 1995, 1890, 1708, 1104, 1263, 1696, 482, 1025, 818, 1619, 1264, 1065, 1930, 1128, 524, 643, 1933, 953, 276, 1101, 1053, 1303, 1010, 1047, 209, 383, 491, 215, 492, 1164, 30, 813, 1392, 770, 341, 1945, 1935, 776, 869, 1973, 189, 2025, 1422, 1626, 1184, 1103, 4, 1905, 1288, 1832, 1977, 1004, 1604, 614, 532, 769, 1609, 1528, 829, 1505, 490, 1638, 1656, 1270, 1717, 374, 316, 862, 1302, 120, 1280, 1599, 1487, 101, 1708, 889, 735, 1662, 1412, 998, 506, 1082, 1391, 1468, 493, 974, 1600, 168, 972, 1989, 1169, 704, 650, 2030, 900, 1285, 51, 1753, 747, 1612, 180, 57, 953, 1215, 252, 127, 280, 780, 1653, 223, 1761, 1220, 568, 1574, 356, 6, 58, 1382, 566, 512, 212, 636, 1621, 270, 1894, 467, 1214, 1350, 1157, 1515, 1325, 1893, 1135, 568, 1970, 296, 1781, 900, 1952, 297, 541, 887, 1636, 424, 767, 1443, 945, 1560, 574, 1145, 0)
   );
end process;   
   
end a1;