library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
use ieee.numeric_std.all;
use IEEE.math_real.all;


package XEf_constants_P5_5d is  

type RTab is array(natural range<>) of std_logic_vector(63 downto 0);
type BitTab is array(natural range<>) of std_logic_vector(7 downto 0);

type ff is array(0 to 255, 0 to 10) of integer; -- fixerr fix
type fu is array(0 to 233, 0 to 4) of integer;  -- fixerr unpack
type cp is array(0 to 233, 0 to 5) of integer; 	-- compute pack
type cr is array(0 to 31, 0 to 8) of integer; 	-- compue reduce poly


constant XEf_fixerr_unpack :=
(
(0, 0, 16, 32, 0),
(0, 1, 16, 32, 1),
(0, 2, 16, 32, 2),
(0, 3, 16, 32, 3),
(0, 4, 16, 32, 4),
(0, 5, 16, 32, 5),
(0, 6, 16, 32, 6),
(0, 7, 16, 32, 7),
(0, 8, 16, 33, 0),
(0, 9, 16, 33, 1),
(0, 10, 16, 33, 2),
(0, 11, 16, 33, 3),
(0, 12, 16, 33, 4),
(0, 13, 16, 33, 5),
(0, 14, 16, 33, 6),
(0, 15, 16, 33, 7),
(1, 0, 16, 34, 0),
(1, 1, 16, 34, 1),
(1, 2, 16, 34, 2),
(1, 3, 16, 34, 3),
(1, 4, 16, 34, 4),
(1, 5, 16, 34, 5),
(1, 6, 16, 34, 6),
(1, 7, 16, 34, 7),
(1, 8, 16, 35, 0),
(1, 9, 16, 35, 1),
(1, 10, 16, 35, 2),
(1, 11, 16, 35, 3),
(1, 12, 16, 35, 4),
(1, 13, 16, 35, 5),
(1, 14, 16, 35, 6),
(1, 15, 16, 35, 7),
(2, 0, 17, 36, 0),
(2, 1, 17, 36, 1),
(2, 2, 17, 36, 2),
(2, 3, 17, 36, 3),
(2, 4, 17, 36, 4),
(2, 5, 17, 36, 5),
(2, 6, 17, 36, 6),
(2, 7, 17, 36, 7),
(2, 8, 17, 37, 0),
(2, 9, 17, 37, 1),
(2, 10, 17, 37, 2),
(2, 11, 17, 37, 3),
(2, 12, 17, 37, 4),
(2, 13, 17, 37, 5),
(2, 14, 17, 37, 6),
(2, 15, 17, 37, 7),
(2, 16, 17, 38, 0),
(3, 0, 19, 38, 1),
(3, 1, 19, 38, 2),
(3, 2, 19, 38, 3),
(3, 3, 19, 38, 4),
(3, 4, 19, 38, 5),
(3, 5, 19, 38, 6),
(3, 6, 19, 38, 7),
(3, 7, 19, 39, 0),
(3, 8, 19, 39, 1),
(3, 9, 19, 39, 2),
(3, 10, 19, 39, 3),
(3, 11, 19, 39, 4),
(3, 12, 19, 39, 5),
(3, 13, 19, 39, 6),
(3, 14, 19, 39, 7),
(3, 15, 19, 40, 0),
(3, 16, 19, 40, 1),
(3, 17, 19, 40, 2),
(3, 18, 19, 40, 3),
(4, 0, 21, 40, 4),
(4, 1, 21, 40, 5),
(4, 2, 21, 40, 6),
(4, 3, 21, 40, 7),
(4, 4, 21, 41, 0),
(4, 5, 21, 41, 1),
(4, 6, 21, 41, 2),
(4, 7, 21, 41, 3),
(4, 8, 21, 41, 4),
(4, 9, 21, 41, 5),
(4, 10, 21, 41, 6),
(4, 11, 21, 41, 7),
(4, 12, 21, 42, 0),
(4, 13, 21, 42, 1),
(4, 14, 21, 42, 2),
(4, 15, 21, 42, 3),
(4, 16, 21, 42, 4),
(4, 17, 21, 42, 5),
(4, 18, 21, 42, 6),
(4, 19, 21, 42, 7),
(4, 20, 21, 43, 0),
(5, 0, 23, 43, 1),
(5, 1, 23, 43, 2),
(5, 2, 23, 43, 3),
(5, 3, 23, 43, 4),
(5, 4, 23, 43, 5),
(5, 5, 23, 43, 6),
(5, 6, 23, 43, 7),
(5, 7, 23, 44, 0),
(5, 8, 23, 44, 1),
(5, 9, 23, 44, 2),
(5, 10, 23, 44, 3),
(5, 11, 23, 44, 4),
(5, 12, 23, 44, 5),
(5, 13, 23, 44, 6),
(5, 14, 23, 44, 7),
(5, 15, 23, 45, 0),
(5, 16, 23, 45, 1),
(5, 17, 23, 45, 2),
(5, 18, 23, 45, 3),
(5, 19, 23, 45, 4),
(5, 20, 23, 45, 5),
(5, 21, 23, 45, 6),
(5, 22, 23, 45, 7),
(6, 0, 25, 46, 0),
(6, 1, 25, 46, 1),
(6, 2, 25, 46, 2),
(6, 3, 25, 46, 3),
(6, 4, 25, 46, 4),
(6, 5, 25, 46, 5),
(6, 6, 25, 46, 6),
(6, 7, 25, 46, 7),
(6, 8, 25, 47, 0),
(6, 9, 25, 47, 1),
(6, 10, 25, 47, 2),
(6, 11, 25, 47, 3),
(6, 12, 25, 47, 4),
(6, 13, 25, 47, 5),
(6, 14, 25, 47, 6),
(6, 15, 25, 47, 7),
(6, 16, 25, 48, 0),
(6, 17, 25, 48, 1),
(6, 18, 25, 48, 2),
(6, 19, 25, 48, 3),
(6, 20, 25, 48, 4),
(6, 21, 25, 48, 5),
(6, 22, 25, 48, 6),
(6, 23, 25, 48, 7),
(6, 24, 25, 49, 0),
(7, 0, 29, 49, 1),
(7, 1, 29, 49, 2),
(7, 2, 29, 49, 3),
(7, 3, 29, 49, 4),
(7, 4, 29, 49, 5),
(7, 5, 29, 49, 6),
(7, 6, 29, 49, 7),
(7, 7, 29, 50, 0),
(7, 8, 29, 50, 1),
(7, 9, 29, 50, 2),
(7, 10, 29, 50, 3),
(7, 11, 29, 50, 4),
(7, 12, 29, 50, 5),
(7, 13, 29, 50, 6),
(7, 14, 29, 50, 7),
(7, 15, 29, 51, 0),
(7, 16, 29, 51, 1),
(7, 17, 29, 51, 2),
(7, 18, 29, 51, 3),
(7, 19, 29, 51, 4),
(7, 20, 29, 51, 5),
(7, 21, 29, 51, 6),
(7, 22, 29, 51, 7),
(7, 23, 29, 52, 0),
(7, 24, 29, 52, 1),
(7, 25, 29, 52, 2),
(7, 26, 29, 52, 3),
(7, 27, 29, 52, 4),
(7, 28, 29, 52, 5),
(8, 0, 31, 52, 6),
(8, 1, 31, 52, 7),
(8, 2, 31, 53, 0),
(8, 3, 31, 53, 1),
(8, 4, 31, 53, 2),
(8, 5, 31, 53, 3),
(8, 6, 31, 53, 4),
(8, 7, 31, 53, 5),
(8, 8, 31, 53, 6),
(8, 9, 31, 53, 7),
(8, 10, 31, 54, 0),
(8, 11, 31, 54, 1),
(8, 12, 31, 54, 2),
(8, 13, 31, 54, 3),
(8, 14, 31, 54, 4),
(8, 15, 31, 54, 5),
(8, 16, 31, 54, 6),
(8, 17, 31, 54, 7),
(8, 18, 31, 55, 0),
(8, 19, 31, 55, 1),
(8, 20, 31, 55, 2),
(8, 21, 31, 55, 3),
(8, 22, 31, 55, 4),
(8, 23, 31, 55, 5),
(8, 24, 31, 55, 6),
(8, 25, 31, 55, 7),
(8, 26, 31, 56, 0),
(8, 27, 31, 56, 1),
(8, 28, 31, 56, 2),
(8, 29, 31, 56, 3),
(8, 30, 31, 56, 4),
(9, 0, 37, 56, 5),
(9, 1, 37, 56, 6),
(9, 2, 37, 56, 7),
(9, 3, 37, 57, 0),
(9, 4, 37, 57, 1),
(9, 5, 37, 57, 2),
(9, 6, 37, 57, 3),
(9, 7, 37, 57, 4),
(9, 8, 37, 57, 5),
(9, 9, 37, 57, 6),
(9, 10, 37, 57, 7),
(9, 11, 37, 58, 0),
(9, 12, 37, 58, 1),
(9, 13, 37, 58, 2),
(9, 14, 37, 58, 3),
(9, 15, 37, 58, 4),
(9, 16, 37, 58, 5),
(9, 17, 37, 58, 6),
(9, 18, 37, 58, 7),
(9, 19, 37, 59, 0),
(9, 20, 37, 59, 1),
(9, 21, 37, 59, 2),
(9, 22, 37, 59, 3),
(9, 23, 37, 59, 4),
(9, 24, 37, 59, 5),
(9, 25, 37, 59, 6),
(9, 26, 37, 59, 7),
(9, 27, 37, 60, 0),
(9, 28, 37, 60, 1),
(9, 29, 37, 60, 2),
(9, 30, 37, 60, 3),
(9, 31, 37, 60, 4),
(9, 32, 37, 60, 5),
(9, 33, 37, 60, 6),
(9, 34, 37, 60, 7),
(9, 35, 37, 61, 0),
(9, 36, 37, 61, 1)
);


constant XEf_fixerr_tab : ff :=
(
( 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0), 
( 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1), 
( 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 2), 
( 0, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 3), 
( 0, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4), 
( 0, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5), 
( 0, 6, 6, 6, 6, 6, 6, 6, 6, 6, 0, 6), 
( 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 7), 
( 0, 8, 8, 8, 8, 8, 8, 8, 8, 8, 1, 0), 
( 0, 9, 9, 9, 9, 9, 9, 9, 9, 9, 1, 1), 
( 0, 10, 10, 10, 10, 10, 10, 10, 10, 10, 1, 2), 
( 0, 11, 11, 11, 11, 11, 11, 11, 11, 11, 1, 3), 
( 0, 12, 12, 12, 12, 12, 12, 12, 12, 12, 1, 4), 
( 0, 13, 13, 13, 13, 13, 13, 13, 13, 13, 1, 5), 
( 0, 14, 14, 14, 14, 14, 14, 14, 14, 14, 1, 6), 
( 0, 15, 15, 15, 15, 15, 15, 15, 15, 15, 1, 7), 
( 1, 0, 16, 16, 16, 16, 16, 16, 16, 16, 2, 0), 
( 1, 1, 0, 17, 17, 17, 17, 17, 17, 17, 2, 1), 
( 1, 2, 1, 18, 18, 18, 18, 18, 18, 18, 2, 2), 
( 1, 3, 2, 0, 19, 19, 19, 19, 19, 19, 2, 3), 
( 1, 4, 3, 1, 20, 20, 20, 20, 20, 20, 2, 4), 
( 1, 5, 4, 2, 0, 21, 21, 21, 21, 21, 2, 5), 
( 1, 6, 5, 3, 1, 22, 22, 22, 22, 22, 2, 6), 
( 1, 7, 6, 4, 2, 0, 23, 23, 23, 23, 2, 7), 
( 1, 8, 7, 5, 3, 1, 24, 24, 24, 24, 3, 0), 
( 1, 9, 8, 6, 4, 2, 0, 25, 25, 25, 3, 1), 
( 1, 10, 9, 7, 5, 3, 1, 26, 26, 26, 3, 2), 
( 1, 11, 10, 8, 6, 4, 2, 27, 27, 27, 3, 3), 
( 1, 12, 11, 9, 7, 5, 3, 28, 28, 28, 3, 4), 
( 1, 13, 12, 10, 8, 6, 4, 0, 29, 29, 3, 5), 
( 1, 14, 13, 11, 9, 7, 5, 1, 30, 30, 3, 6), 
( 1, 15, 14, 12, 10, 8, 6, 2, 0, 31, 3, 7), 
( 2, 0, 15, 13, 11, 9, 7, 3, 1, 32, 4, 0), 
( 2, 1, 16, 14, 12, 10, 8, 4, 2, 33, 4, 1), 
( 2, 2, 0, 15, 13, 11, 9, 5, 3, 34, 4, 2), 
( 2, 3, 1, 16, 14, 12, 10, 6, 4, 35, 4, 3), 
( 2, 4, 2, 17, 15, 13, 11, 7, 5, 36, 4, 4), 
( 2, 5, 3, 18, 16, 14, 12, 8, 6, 0, 4, 5), 
( 2, 6, 4, 0, 17, 15, 13, 9, 7, 1, 4, 6), 
( 2, 7, 5, 1, 18, 16, 14, 10, 8, 2, 4, 7), 
( 2, 8, 6, 2, 19, 17, 15, 11, 9, 3, 5, 0), 
( 2, 9, 7, 3, 20, 18, 16, 12, 10, 4, 5, 1), 
( 2, 10, 8, 4, 0, 19, 17, 13, 11, 5, 5, 2), 
( 2, 11, 9, 5, 1, 20, 18, 14, 12, 6, 5, 3), 
( 2, 12, 10, 6, 2, 21, 19, 15, 13, 7, 5, 4), 
( 2, 13, 11, 7, 3, 22, 20, 16, 14, 8, 5, 5), 
( 2, 14, 12, 8, 4, 0, 21, 17, 15, 9, 5, 6), 
( 2, 15, 13, 9, 5, 1, 22, 18, 16, 10, 5, 7), 
( 3, 0, 14, 10, 6, 2, 23, 19, 17, 11, 6, 0), 
( 3, 1, 15, 11, 7, 3, 24, 20, 18, 12, 6, 1), 
( 3, 2, 16, 12, 8, 4, 0, 21, 19, 13, 6, 2), 
( 3, 3, 0, 13, 9, 5, 1, 22, 20, 14, 6, 3), 
( 3, 4, 1, 14, 10, 6, 2, 23, 21, 15, 6, 4), 
( 3, 5, 2, 15, 11, 7, 3, 24, 22, 16, 6, 5), 
( 3, 6, 3, 16, 12, 8, 4, 25, 23, 17, 6, 6), 
( 3, 7, 4, 17, 13, 9, 5, 26, 24, 18, 6, 7), 
( 3, 8, 5, 18, 14, 10, 6, 27, 25, 19, 7, 0), 
( 3, 9, 6, 0, 15, 11, 7, 28, 26, 20, 7, 1), 
( 3, 10, 7, 1, 16, 12, 8, 0, 27, 21, 7, 2), 
( 3, 11, 8, 2, 17, 13, 9, 1, 28, 22, 7, 3), 
( 3, 12, 9, 3, 18, 14, 10, 2, 29, 23, 7, 4), 
( 3, 13, 10, 4, 19, 15, 11, 3, 30, 24, 7, 5), 
( 3, 14, 11, 5, 20, 16, 12, 4, 0, 25, 7, 6), 
( 3, 15, 12, 6, 0, 17, 13, 5, 1, 26, 7, 7), 
( 4, 0, 13, 7, 1, 18, 14, 6, 2, 27, 8, 0), 
( 4, 1, 14, 8, 2, 19, 15, 7, 3, 28, 8, 1), 
( 4, 2, 15, 9, 3, 20, 16, 8, 4, 29, 8, 2), 
( 4, 3, 16, 10, 4, 21, 17, 9, 5, 30, 8, 3), 
( 4, 4, 0, 11, 5, 22, 18, 10, 6, 31, 8, 4), 
( 4, 5, 1, 12, 6, 0, 19, 11, 7, 32, 8, 5), 
( 4, 6, 2, 13, 7, 1, 20, 12, 8, 33, 8, 6), 
( 4, 7, 3, 14, 8, 2, 21, 13, 9, 34, 8, 7), 
( 4, 8, 4, 15, 9, 3, 22, 14, 10, 35, 9, 0), 
( 4, 9, 5, 16, 10, 4, 23, 15, 11, 36, 9, 1), 
( 4, 10, 6, 17, 11, 5, 24, 16, 12, 0, 9, 2), 
( 4, 11, 7, 18, 12, 6, 0, 17, 13, 1, 9, 3), 
( 4, 12, 8, 0, 13, 7, 1, 18, 14, 2, 9, 4), 
( 4, 13, 9, 1, 14, 8, 2, 19, 15, 3, 9, 5), 
( 4, 14, 10, 2, 15, 9, 3, 20, 16, 4, 9, 6), 
( 4, 15, 11, 3, 16, 10, 4, 21, 17, 5, 9, 7), 
( 5, 0, 12, 4, 17, 11, 5, 22, 18, 6, 10, 0), 
( 5, 1, 13, 5, 18, 12, 6, 23, 19, 7, 10, 1), 
( 5, 2, 14, 6, 19, 13, 7, 24, 20, 8, 10, 2), 
( 5, 3, 15, 7, 20, 14, 8, 25, 21, 9, 10, 3), 
( 5, 4, 16, 8, 0, 15, 9, 26, 22, 10, 10, 4), 
( 5, 5, 0, 9, 1, 16, 10, 27, 23, 11, 10, 5), 
( 5, 6, 1, 10, 2, 17, 11, 28, 24, 12, 10, 6), 
( 5, 7, 2, 11, 3, 18, 12, 0, 25, 13, 10, 7), 
( 5, 8, 3, 12, 4, 19, 13, 1, 26, 14, 11, 0), 
( 5, 9, 4, 13, 5, 20, 14, 2, 27, 15, 11, 1), 
( 5, 10, 5, 14, 6, 21, 15, 3, 28, 16, 11, 2), 
( 5, 11, 6, 15, 7, 22, 16, 4, 29, 17, 11, 3), 
( 5, 12, 7, 16, 8, 0, 17, 5, 30, 18, 11, 4), 
( 5, 13, 8, 17, 9, 1, 18, 6, 0, 19, 11, 5), 
( 5, 14, 9, 18, 10, 2, 19, 7, 1, 20, 11, 6), 
( 5, 15, 10, 0, 11, 3, 20, 8, 2, 21, 11, 7), 
( 6, 0, 11, 1, 12, 4, 21, 9, 3, 22, 12, 0), 
( 6, 1, 12, 2, 13, 5, 22, 10, 4, 23, 12, 1), 
( 6, 2, 13, 3, 14, 6, 23, 11, 5, 24, 12, 2), 
( 6, 3, 14, 4, 15, 7, 24, 12, 6, 25, 12, 3), 
( 6, 4, 15, 5, 16, 8, 0, 13, 7, 26, 12, 4), 
( 6, 5, 16, 6, 17, 9, 1, 14, 8, 27, 12, 5), 
( 6, 6, 0, 7, 18, 10, 2, 15, 9, 28, 12, 6), 
( 6, 7, 1, 8, 19, 11, 3, 16, 10, 29, 12, 7), 
( 6, 8, 2, 9, 20, 12, 4, 17, 11, 30, 13, 0), 
( 6, 9, 3, 10, 0, 13, 5, 18, 12, 31, 13, 1), 
( 6, 10, 4, 11, 1, 14, 6, 19, 13, 32, 13, 2), 
( 6, 11, 5, 12, 2, 15, 7, 20, 14, 33, 13, 3), 
( 6, 12, 6, 13, 3, 16, 8, 21, 15, 34, 13, 4), 
( 6, 13, 7, 14, 4, 17, 9, 22, 16, 35, 13, 5), 
( 6, 14, 8, 15, 5, 18, 10, 23, 17, 36, 13, 6), 
( 6, 15, 9, 16, 6, 19, 11, 24, 18, 0, 13, 7), 
( 7, 0, 10, 17, 7, 20, 12, 25, 19, 1, 14, 0), 
( 7, 1, 11, 18, 8, 21, 13, 26, 20, 2, 14, 1), 
( 7, 2, 12, 0, 9, 22, 14, 27, 21, 3, 14, 2), 
( 7, 3, 13, 1, 10, 0, 15, 28, 22, 4, 14, 3), 
( 7, 4, 14, 2, 11, 1, 16, 0, 23, 5, 14, 4), 
( 7, 5, 15, 3, 12, 2, 17, 1, 24, 6, 14, 5), 
( 7, 6, 16, 4, 13, 3, 18, 2, 25, 7, 14, 6), 
( 7, 7, 0, 5, 14, 4, 19, 3, 26, 8, 14, 7), 
( 7, 8, 1, 6, 15, 5, 20, 4, 27, 9, 15, 0), 
( 7, 9, 2, 7, 16, 6, 21, 5, 28, 10, 15, 1), 
( 7, 10, 3, 8, 17, 7, 22, 6, 29, 11, 15, 2), 
( 7, 11, 4, 9, 18, 8, 23, 7, 30, 12, 15, 3), 
( 7, 12, 5, 10, 19, 9, 24, 8, 0, 13, 15, 4), 
( 7, 13, 6, 11, 20, 10, 0, 9, 1, 14, 15, 5), 
( 7, 14, 7, 12, 0, 11, 1, 10, 2, 15, 15, 6), 
( 7, 15, 8, 13, 1, 12, 2, 11, 3, 16, 15, 7), 
( 8, 0, 9, 14, 2, 13, 3, 12, 4, 17, 16, 0), 
( 8, 1, 10, 15, 3, 14, 4, 13, 5, 18, 16, 1), 
( 8, 2, 11, 16, 4, 15, 5, 14, 6, 19, 16, 2), 
( 8, 3, 12, 17, 5, 16, 6, 15, 7, 20, 16, 3), 
( 8, 4, 13, 18, 6, 17, 7, 16, 8, 21, 16, 4), 
( 8, 5, 14, 0, 7, 18, 8, 17, 9, 22, 16, 5), 
( 8, 6, 15, 1, 8, 19, 9, 18, 10, 23, 16, 6), 
( 8, 7, 16, 2, 9, 20, 10, 19, 11, 24, 16, 7), 
( 8, 8, 0, 3, 10, 21, 11, 20, 12, 25, 17, 0), 
( 8, 9, 1, 4, 11, 22, 12, 21, 13, 26, 17, 1), 
( 8, 10, 2, 5, 12, 0, 13, 22, 14, 27, 17, 2), 
( 8, 11, 3, 6, 13, 1, 14, 23, 15, 28, 17, 3), 
( 8, 12, 4, 7, 14, 2, 15, 24, 16, 29, 17, 4), 
( 8, 13, 5, 8, 15, 3, 16, 25, 17, 30, 17, 5), 
( 8, 14, 6, 9, 16, 4, 17, 26, 18, 31, 17, 6), 
( 8, 15, 7, 10, 17, 5, 18, 27, 19, 32, 17, 7), 
( 9, 0, 8, 11, 18, 6, 19, 28, 20, 33, 18, 0), 
( 9, 1, 9, 12, 19, 7, 20, 0, 21, 34, 18, 1), 
( 9, 2, 10, 13, 20, 8, 21, 1, 22, 35, 18, 2), 
( 9, 3, 11, 14, 0, 9, 22, 2, 23, 36, 18, 3), 
( 9, 4, 12, 15, 1, 10, 23, 3, 24, 0, 18, 4), 
( 9, 5, 13, 16, 2, 11, 24, 4, 25, 1, 18, 5), 
( 9, 6, 14, 17, 3, 12, 0, 5, 26, 2, 18, 6), 
( 9, 7, 15, 18, 4, 13, 1, 6, 27, 3, 18, 7), 
( 9, 8, 16, 0, 5, 14, 2, 7, 28, 4, 19, 0), 
( 9, 9, 0, 1, 6, 15, 3, 8, 29, 5, 19, 1), 
( 9, 10, 1, 2, 7, 16, 4, 9, 30, 6, 19, 2), 
( 9, 11, 2, 3, 8, 17, 5, 10, 0, 7, 19, 3), 
( 9, 12, 3, 4, 9, 18, 6, 11, 1, 8, 19, 4), 
( 9, 13, 4, 5, 10, 19, 7, 12, 2, 9, 19, 5), 
( 9, 14, 5, 6, 11, 20, 8, 13, 3, 10, 19, 6), 
( 9, 15, 6, 7, 12, 21, 9, 14, 4, 11, 19, 7), 
( 10, 0, 7, 8, 13, 22, 10, 15, 5, 12, 20, 0), 
( 10, 1, 8, 9, 14, 0, 11, 16, 6, 13, 20, 1), 
( 10, 2, 9, 10, 15, 1, 12, 17, 7, 14, 20, 2), 
( 10, 3, 10, 11, 16, 2, 13, 18, 8, 15, 20, 3), 
( 10, 4, 11, 12, 17, 3, 14, 19, 9, 16, 20, 4), 
( 10, 5, 12, 13, 18, 4, 15, 20, 10, 17, 20, 5), 
( 10, 6, 13, 14, 19, 5, 16, 21, 11, 18, 20, 6), 
( 10, 7, 14, 15, 20, 6, 17, 22, 12, 19, 20, 7), 
( 10, 8, 15, 16, 0, 7, 18, 23, 13, 20, 21, 0), 
( 10, 9, 16, 17, 1, 8, 19, 24, 14, 21, 21, 1), 
( 10, 10, 0, 18, 2, 9, 20, 25, 15, 22, 21, 2), 
( 10, 11, 1, 0, 3, 10, 21, 26, 16, 23, 21, 3), 
( 10, 12, 2, 1, 4, 11, 22, 27, 17, 24, 21, 4), 
( 10, 13, 3, 2, 5, 12, 23, 28, 18, 25, 21, 5), 
( 10, 14, 4, 3, 6, 13, 24, 0, 19, 26, 21, 6), 
( 10, 15, 5, 4, 7, 14, 0, 1, 20, 27, 21, 7), 
( 11, 0, 6, 5, 8, 15, 1, 2, 21, 28, 22, 0), 
( 11, 1, 7, 6, 9, 16, 2, 3, 22, 29, 22, 1), 
( 11, 2, 8, 7, 10, 17, 3, 4, 23, 30, 22, 2), 
( 11, 3, 9, 8, 11, 18, 4, 5, 24, 31, 22, 3), 
( 11, 4, 10, 9, 12, 19, 5, 6, 25, 32, 22, 4), 
( 11, 5, 11, 10, 13, 20, 6, 7, 26, 33, 22, 5), 
( 11, 6, 12, 11, 14, 21, 7, 8, 27, 34, 22, 6), 
( 11, 7, 13, 12, 15, 22, 8, 9, 28, 35, 22, 7), 
( 11, 8, 14, 13, 16, 0, 9, 10, 29, 36, 23, 0), 
( 11, 9, 15, 14, 17, 1, 10, 11, 30, 0, 23, 1), 
( 11, 10, 16, 15, 18, 2, 11, 12, 0, 1, 23, 2), 
( 11, 11, 0, 16, 19, 3, 12, 13, 1, 2, 23, 3), 
( 11, 12, 1, 17, 20, 4, 13, 14, 2, 3, 23, 4), 
( 11, 13, 2, 18, 0, 5, 14, 15, 3, 4, 23, 5), 
( 11, 14, 3, 0, 1, 6, 15, 16, 4, 5, 23, 6), 
( 11, 15, 4, 1, 2, 7, 16, 17, 5, 6, 23, 7), 
( 12, 0, 5, 2, 3, 8, 17, 18, 6, 7, 24, 0), 
( 12, 1, 6, 3, 4, 9, 18, 19, 7, 8, 24, 1), 
( 12, 2, 7, 4, 5, 10, 19, 20, 8, 9, 24, 2), 
( 12, 3, 8, 5, 6, 11, 20, 21, 9, 10, 24, 3), 
( 12, 4, 9, 6, 7, 12, 21, 22, 10, 11, 24, 4), 
( 12, 5, 10, 7, 8, 13, 22, 23, 11, 12, 24, 5), 
( 12, 6, 11, 8, 9, 14, 23, 24, 12, 13, 24, 6), 
( 12, 7, 12, 9, 10, 15, 24, 25, 13, 14, 24, 7), 
( 12, 8, 13, 10, 11, 16, 0, 26, 14, 15, 25, 0), 
( 12, 9, 14, 11, 12, 17, 1, 27, 15, 16, 25, 1), 
( 12, 10, 15, 12, 13, 18, 2, 28, 16, 17, 25, 2), 
( 12, 11, 16, 13, 14, 19, 3, 0, 17, 18, 25, 3), 
( 12, 12, 0, 14, 15, 20, 4, 1, 18, 19, 25, 4), 
( 12, 13, 1, 15, 16, 21, 5, 2, 19, 20, 25, 5), 
( 12, 14, 2, 16, 17, 22, 6, 3, 20, 21, 25, 6), 
( 12, 15, 3, 17, 18, 0, 7, 4, 21, 22, 25, 7), 
( 13, 0, 4, 18, 19, 1, 8, 5, 22, 23, 26, 0), 
( 13, 1, 5, 0, 20, 2, 9, 6, 23, 24, 26, 1), 
( 13, 2, 6, 1, 0, 3, 10, 7, 24, 25, 26, 2), 
( 13, 3, 7, 2, 1, 4, 11, 8, 25, 26, 26, 3), 
( 13, 4, 8, 3, 2, 5, 12, 9, 26, 27, 26, 4), 
( 13, 5, 9, 4, 3, 6, 13, 10, 27, 28, 26, 5), 
( 13, 6, 10, 5, 4, 7, 14, 11, 28, 29, 26, 6), 
( 13, 7, 11, 6, 5, 8, 15, 12, 29, 30, 26, 7), 
( 13, 8, 12, 7, 6, 9, 16, 13, 30, 31, 27, 0), 
( 13, 9, 13, 8, 7, 10, 17, 14, 0, 32, 27, 1), 
( 13, 10, 14, 9, 8, 11, 18, 15, 1, 33, 27, 2), 
( 13, 11, 15, 10, 9, 12, 19, 16, 2, 34, 27, 3), 
( 13, 12, 16, 11, 10, 13, 20, 17, 3, 35, 27, 4), 
( 13, 13, 0, 12, 11, 14, 21, 18, 4, 36, 27, 5), 
( 13, 14, 1, 13, 12, 15, 22, 19, 5, 0, 27, 6), 
( 13, 15, 2, 14, 13, 16, 23, 20, 6, 1, 27, 7), 
( 14, 0, 3, 15, 14, 17, 24, 21, 7, 2, 28, 0), 
( 14, 1, 4, 16, 15, 18, 0, 22, 8, 3, 28, 1), 
( 14, 2, 5, 17, 16, 19, 1, 23, 9, 4, 28, 2), 
( 14, 3, 6, 18, 17, 20, 2, 24, 10, 5, 28, 3), 
( 14, 4, 7, 0, 18, 21, 3, 25, 11, 6, 28, 4), 
( 14, 5, 8, 1, 19, 22, 4, 26, 12, 7, 28, 5), 
( 14, 6, 9, 2, 20, 0, 5, 27, 13, 8, 28, 6), 
( 14, 7, 10, 3, 0, 1, 6, 28, 14, 9, 28, 7), 
( 14, 8, 11, 4, 1, 2, 7, 0, 15, 10, 29, 0), 
( 14, 9, 12, 5, 2, 3, 8, 1, 16, 11, 29, 1), 
( 14, 10, 13, 6, 3, 4, 9, 2, 17, 12, 29, 2), 
( 14, 11, 14, 7, 4, 5, 10, 3, 18, 13, 29, 3), 
( 14, 12, 15, 8, 5, 6, 11, 4, 19, 14, 29, 4), 
( 14, 13, 16, 9, 6, 7, 12, 5, 20, 15, 29, 5), 
( 14, 14, 0, 10, 7, 8, 13, 6, 21, 16, 29, 6), 
( 14, 15, 1, 11, 8, 9, 14, 7, 22, 17, 29, 7), 
( 15, 0, 2, 12, 9, 10, 15, 8, 23, 18, 30, 0), 
( 15, 1, 3, 13, 10, 11, 16, 9, 24, 19, 30, 1), 
( 15, 2, 4, 14, 11, 12, 17, 10, 25, 20, 30, 2), 
( 15, 3, 5, 15, 12, 13, 18, 11, 26, 21, 30, 3), 
( 15, 4, 6, 16, 13, 14, 19, 12, 27, 22, 30, 4), 
( 15, 5, 7, 17, 14, 15, 20, 13, 28, 23, 30, 5), 
( 15, 6, 8, 18, 15, 16, 21, 14, 29, 24, 30, 6), 
( 15, 7, 9, 0, 16, 17, 22, 15, 30, 25, 30, 7), 
( 15, 8, 10, 1, 17, 18, 23, 16, 0, 26, 31, 0), 
( 15, 9, 11, 2, 18, 19, 24, 17, 1, 27, 31, 1), 
( 15, 10, 12, 3, 19, 20, 0, 18, 2, 28, 31, 2), 
( 15, 11, 13, 4, 20, 21, 1, 19, 3, 29, 31, 3), 
( 15, 12, 14, 5, 0, 22, 2, 20, 4, 30, 31, 4), 
( 15, 13, 15, 6, 1, 0, 3, 21, 5, 31, 31, 5), 
( 15, 14, 16, 7, 2, 1, 4, 22, 6, 32, 31, 6), 
( 15, 15, 0, 8, 3, 2, 5, 23, 7, 33, 31, 7)
);

constant XEf_reduce_poly : cr :=
(
(0, 0, 0, 0, 0, 0, 0, 0, 0),
(8, 8, 8, 8, 8, 8, 8, 8, 8),
(0, 16, 16, 16, 16, 16, 16, 16, 16),
(8, 7, 5, 3, 1, 24, 24, 24, 24),
(0, 15, 13, 11, 9, 7, 3, 1, 32),
(8, 6, 2, 19, 17, 15, 11, 9, 3),
(0, 14, 10, 6, 2, 23, 19, 17, 11),
(8, 5, 18, 14, 10, 6, 27, 25, 19),
(0, 13, 7, 1, 18, 14, 6, 2, 27),
(8, 4, 15, 9, 3, 22, 14, 10, 35),
(0, 12, 4, 17, 11, 5, 22, 18, 6),
(8, 3, 12, 4, 19, 13, 1, 26, 14),
(0, 11, 1, 12, 4, 21, 9, 3, 22),
(8, 2, 9, 20, 12, 4, 17, 11, 30),
(0, 10, 17, 7, 20, 12, 25, 19, 1),
(8, 1, 6, 15, 5, 20, 4, 27, 9),
(0, 9, 14, 2, 13, 3, 12, 4, 17),
(8, 0, 3, 10, 21, 11, 20, 12, 25),
(0, 8, 11, 18, 6, 19, 28, 20, 33),
(8, 16, 0, 5, 14, 2, 7, 28, 4),
(0, 7, 8, 13, 22, 10, 15, 5, 12),
(8, 15, 16, 0, 7, 18, 23, 13, 20),
(0, 6, 5, 8, 15, 1, 2, 21, 28),
(8, 14, 13, 16, 0, 9, 10, 29, 36),
(0, 5, 2, 3, 8, 17, 18, 6, 7),
(8, 13, 10, 11, 16, 0, 26, 14, 15),
(0, 4, 18, 19, 1, 8, 5, 22, 23),
(8, 12, 7, 6, 9, 16, 13, 30, 31),
(0, 3, 15, 14, 17, 24, 21, 7, 2),
(8, 11, 4, 1, 2, 7, 0, 15, 10),
(0, 2, 12, 9, 10, 15, 8, 23, 18),
(8, 10, 1, 17, 18, 23, 16, 0, 26)
);

constant XEf_compute_pack : cp :=
(
(0, 0, 16, 256, 32, 0),
(0, 1, 16, 257, 32, 1),
(0, 2, 16, 258, 32, 2),
(0, 3, 16, 259, 32, 3),
(0, 4, 16, 260, 32, 4),
(0, 5, 16, 261, 32, 5),
(0, 6, 16, 262, 32, 6),
(0, 7, 16, 263, 32, 7),
(0, 8, 16, 264, 33, 0),
(0, 9, 16, 265, 33, 1),
(0, 10, 16, 266, 33, 2),
(0, 11, 16, 267, 33, 3),
(0, 12, 16, 268, 33, 4),
(0, 13, 16, 269, 33, 5),
(0, 14, 16, 270, 33, 6),
(0, 15, 16, 271, 33, 7),
(1, 0, 16, 272, 34, 0),
(1, 1, 16, 273, 34, 1),
(1, 2, 16, 274, 34, 2),
(1, 3, 16, 275, 34, 3),
(1, 4, 16, 276, 34, 4),
(1, 5, 16, 277, 34, 5),
(1, 6, 16, 278, 34, 6),
(1, 7, 16, 279, 34, 7),
(1, 8, 16, 280, 35, 0),
(1, 9, 16, 281, 35, 1),
(1, 10, 16, 282, 35, 2),
(1, 11, 16, 283, 35, 3),
(1, 12, 16, 284, 35, 4),
(1, 13, 16, 285, 35, 5),
(1, 14, 16, 286, 35, 6),
(1, 15, 16, 287, 35, 7),
(2, 0, 17, 288, 36, 0),
(2, 1, 17, 289, 36, 1),
(2, 2, 17, 290, 36, 2),
(2, 3, 17, 291, 36, 3),
(2, 4, 17, 292, 36, 4),
(2, 5, 17, 293, 36, 5),
(2, 6, 17, 294, 36, 6),
(2, 7, 17, 295, 36, 7),
(2, 8, 17, 296, 37, 0),
(2, 9, 17, 297, 37, 1),
(2, 10, 17, 298, 37, 2),
(2, 11, 17, 299, 37, 3),
(2, 12, 17, 300, 37, 4),
(2, 13, 17, 301, 37, 5),
(2, 14, 17, 302, 37, 6),
(2, 15, 17, 303, 37, 7),
(2, 16, 17, 304, 38, 0),
(3, 0, 19, 305, 38, 1),
(3, 1, 19, 306, 38, 2),
(3, 2, 19, 307, 38, 3),
(3, 3, 19, 308, 38, 4),
(3, 4, 19, 309, 38, 5),
(3, 5, 19, 310, 38, 6),
(3, 6, 19, 311, 38, 7),
(3, 7, 19, 312, 39, 0),
(3, 8, 19, 313, 39, 1),
(3, 9, 19, 314, 39, 2),
(3, 10, 19, 315, 39, 3),
(3, 11, 19, 316, 39, 4),
(3, 12, 19, 317, 39, 5),
(3, 13, 19, 318, 39, 6),
(3, 14, 19, 319, 39, 7),
(3, 15, 19, 320, 40, 0),
(3, 16, 19, 321, 40, 1),
(3, 17, 19, 322, 40, 2),
(3, 18, 19, 323, 40, 3),
(4, 0, 21, 324, 40, 4),
(4, 1, 21, 325, 40, 5),
(4, 2, 21, 326, 40, 6),
(4, 3, 21, 327, 40, 7),
(4, 4, 21, 328, 41, 0),
(4, 5, 21, 329, 41, 1),
(4, 6, 21, 330, 41, 2),
(4, 7, 21, 331, 41, 3),
(4, 8, 21, 332, 41, 4),
(4, 9, 21, 333, 41, 5),
(4, 10, 21, 334, 41, 6),
(4, 11, 21, 335, 41, 7),
(4, 12, 21, 336, 42, 0),
(4, 13, 21, 337, 42, 1),
(4, 14, 21, 338, 42, 2),
(4, 15, 21, 339, 42, 3),
(4, 16, 21, 340, 42, 4),
(4, 17, 21, 341, 42, 5),
(4, 18, 21, 342, 42, 6),
(4, 19, 21, 343, 42, 7),
(4, 20, 21, 344, 43, 0),
(5, 0, 23, 345, 43, 1),
(5, 1, 23, 346, 43, 2),
(5, 2, 23, 347, 43, 3),
(5, 3, 23, 348, 43, 4),
(5, 4, 23, 349, 43, 5),
(5, 5, 23, 350, 43, 6),
(5, 6, 23, 351, 43, 7),
(5, 7, 23, 352, 44, 0),
(5, 8, 23, 353, 44, 1),
(5, 9, 23, 354, 44, 2),
(5, 10, 23, 355, 44, 3),
(5, 11, 23, 356, 44, 4),
(5, 12, 23, 357, 44, 5),
(5, 13, 23, 358, 44, 6),
(5, 14, 23, 359, 44, 7),
(5, 15, 23, 360, 45, 0),
(5, 16, 23, 361, 45, 1),
(5, 17, 23, 362, 45, 2),
(5, 18, 23, 363, 45, 3),
(5, 19, 23, 364, 45, 4),
(5, 20, 23, 365, 45, 5),
(5, 21, 23, 366, 45, 6),
(5, 22, 23, 367, 45, 7),
(6, 0, 25, 368, 46, 0),
(6, 1, 25, 369, 46, 1),
(6, 2, 25, 370, 46, 2),
(6, 3, 25, 371, 46, 3),
(6, 4, 25, 372, 46, 4),
(6, 5, 25, 373, 46, 5),
(6, 6, 25, 374, 46, 6),
(6, 7, 25, 375, 46, 7),
(6, 8, 25, 376, 47, 0),
(6, 9, 25, 377, 47, 1),
(6, 10, 25, 378, 47, 2),
(6, 11, 25, 379, 47, 3),
(6, 12, 25, 380, 47, 4),
(6, 13, 25, 381, 47, 5),
(6, 14, 25, 382, 47, 6),
(6, 15, 25, 383, 47, 7),
(6, 16, 25, 384, 48, 0),
(6, 17, 25, 385, 48, 1),
(6, 18, 25, 386, 48, 2),
(6, 19, 25, 387, 48, 3),
(6, 20, 25, 388, 48, 4),
(6, 21, 25, 389, 48, 5),
(6, 22, 25, 390, 48, 6),
(6, 23, 25, 391, 48, 7),
(6, 24, 25, 392, 49, 0),
(7, 0, 29, 393, 49, 1),
(7, 1, 29, 394, 49, 2),
(7, 2, 29, 395, 49, 3),
(7, 3, 29, 396, 49, 4),
(7, 4, 29, 397, 49, 5),
(7, 5, 29, 398, 49, 6),
(7, 6, 29, 399, 49, 7),
(7, 7, 29, 400, 50, 0),
(7, 8, 29, 401, 50, 1),
(7, 9, 29, 402, 50, 2),
(7, 10, 29, 403, 50, 3),
(7, 11, 29, 404, 50, 4),
(7, 12, 29, 405, 50, 5),
(7, 13, 29, 406, 50, 6),
(7, 14, 29, 407, 50, 7),
(7, 15, 29, 408, 51, 0),
(7, 16, 29, 409, 51, 1),
(7, 17, 29, 410, 51, 2),
(7, 18, 29, 411, 51, 3),
(7, 19, 29, 412, 51, 4),
(7, 20, 29, 413, 51, 5),
(7, 21, 29, 414, 51, 6),
(7, 22, 29, 415, 51, 7),
(7, 23, 29, 416, 52, 0),
(7, 24, 29, 417, 52, 1),
(7, 25, 29, 418, 52, 2),
(7, 26, 29, 419, 52, 3),
(7, 27, 29, 420, 52, 4),
(7, 28, 29, 421, 52, 5),
(8, 0, 31, 422, 52, 6),
(8, 1, 31, 423, 52, 7),
(8, 2, 31, 424, 53, 0),
(8, 3, 31, 425, 53, 1),
(8, 4, 31, 426, 53, 2),
(8, 5, 31, 427, 53, 3),
(8, 6, 31, 428, 53, 4),
(8, 7, 31, 429, 53, 5),
(8, 8, 31, 430, 53, 6),
(8, 9, 31, 431, 53, 7),
(8, 10, 31, 432, 54, 0),
(8, 11, 31, 433, 54, 1),
(8, 12, 31, 434, 54, 2),
(8, 13, 31, 435, 54, 3),
(8, 14, 31, 436, 54, 4),
(8, 15, 31, 437, 54, 5),
(8, 16, 31, 438, 54, 6),
(8, 17, 31, 439, 54, 7),
(8, 18, 31, 440, 55, 0),
(8, 19, 31, 441, 55, 1),
(8, 20, 31, 442, 55, 2),
(8, 21, 31, 443, 55, 3),
(8, 22, 31, 444, 55, 4),
(8, 23, 31, 445, 55, 5),
(8, 24, 31, 446, 55, 6),
(8, 25, 31, 447, 55, 7),
(8, 26, 31, 448, 56, 0),
(8, 27, 31, 449, 56, 1),
(8, 28, 31, 450, 56, 2),
(8, 29, 31, 451, 56, 3),
(8, 30, 31, 452, 56, 4),
(9, 0, 37, 453, 56, 5),
(9, 1, 37, 454, 56, 6),
(9, 2, 37, 455, 56, 7),
(9, 3, 37, 456, 57, 0),
(9, 4, 37, 457, 57, 1),
(9, 5, 37, 458, 57, 2),
(9, 6, 37, 459, 57, 3),
(9, 7, 37, 460, 57, 4),
(9, 8, 37, 461, 57, 5),
(9, 9, 37, 462, 57, 6),
(9, 10, 37, 463, 57, 7),
(9, 11, 37, 464, 58, 0),
(9, 12, 37, 465, 58, 1),
(9, 13, 37, 466, 58, 2),
(9, 14, 37, 467, 58, 3),
(9, 15, 37, 468, 58, 4),
(9, 16, 37, 469, 58, 5),
(9, 17, 37, 470, 58, 6),
(9, 18, 37, 471, 58, 7),
(9, 19, 37, 472, 59, 0),
(9, 20, 37, 473, 59, 1),
(9, 21, 37, 474, 59, 2),
(9, 22, 37, 475, 59, 3),
(9, 23, 37, 476, 59, 4),
(9, 24, 37, 477, 59, 5),
(9, 25, 37, 478, 59, 6),
(9, 26, 37, 479, 59, 7),
(9, 27, 37, 480, 60, 0),
(9, 28, 37, 481, 60, 1),
(9, 29, 37, 482, 60, 2),
(9, 30, 37, 483, 60, 3),
(9, 31, 37, 484, 60, 4),
(9, 32, 37, 485, 60, 5),
(9, 33, 37, 486, 60, 6),
(9, 34, 37, 487, 60, 7),
(9, 35, 37, 488, 61, 0),
(9, 36, 37, 489, 61, 1)
);







end package;
