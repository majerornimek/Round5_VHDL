library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
use ieee.numeric_std.all;

library work;
use work.Round5_constants.all;

entity Mul_Poly_TB is
end entity; 

architecture a1 of Mul_Poly_TB is 
component Mul_Poly is 
	port (
		PolyA	: in NTRUPoly(PolyDegree downto 0);
		PolyB	: in Trinomial(PolyDegree downto 0); 
		clk		: in std_logic;
		Start	: in std_logic;
		Rst		: in std_logic;
		OpType	: in std_logic;
		Done	: out std_logic;
		LongRes	: out NTRUPoly(PolyDegree downto 0);
		ShortRes: out ShortPoly(PolyDegree downto 0)
	);
end component;
signal inA, outC : NTRUPoly(PolyDegree downto 0);
signal inB : Trinomial(PolyDegree downto  0); 
signal outS : ShortPoly(PolyDegree downto  0);
signal clk, start_tmp, rst_tmp, op_tmp, done_tmp : std_logic;
constant CLK_PERIOD : time := 10 ps;
type input_array is array(PolyDegree downto 0) of integer;

begin

 clk_process :process
   begin
        clk <= '0';
        wait for CLK_PERIOD/2;  --for half of clock period clk stays at '0'.
        clk <= '1';
        wait for CLK_PERIOD/2;  --for next half of clock period clk stays at '1'.
   end process;
   
   uut: Mul_Poly port map(
    	PolyA	=> inA,
		PolyB	=> inB,
		clk		=> clk,
		Start	=> start_tmp,
		Rst		=> rst_tmp,
		OpType	=> op_tmp,
		Done	=> done_tmp,
		LongRes	=> outC,
		ShortRes=> outS
   );
   
process
	
	procedure check_poly_mul( 	constant PolyA	: in input_array; -- v1
								constant PolyB 	: in input_array; -- v2
								constant typ	: in std_logic; -- norm of v1
								constant res_ex	: in input_array) is
		variable res: input_array;
	begin
		GG: for i in PolyDegree downto 0 loop
			inA(i) <= std_logic_vector(to_signed(PolyA(i), LongModLen));
			inB(i) <= std_logic_vector(to_signed(PolyB(i), 2));
		end loop GG;
		
		wait for CLK_PERIOD;
		rst_tmp <= '1';
		op_tmp <= typ;
		wait for CLK_PERIOD;
		rst_tmp <= '0';
		start_tmp <= '1';
		wait for CLK_PERIOD*700;
		start_tmp <= '0';
		wait for CLK_PERIOD;
		
--		RR: for i in NUM_OF_ELEMENTS-1 downto 0 loop
--			res(i) = to_integer(signed(outC(i)));
--		end loop RR;
--		assert res = res_ex
--		report 	"Unexpected result: " --&
----				"IN1 = " & integer'image(in1) & "; " &
----				"IN2 = " & integer'image(in2) & "; " &
----				"MUL = " & integer'image(res) & "; " &
----				"MUL_expected = " & integer'image(res_ex)
--		severity error;
	end procedure check_poly_mul;
	
	
begin
	

    --618
   check_poly_mul((1400,7,1894,1015,591,475,489,1030,805,1023,1725,1419,277,492,1599,1959,423,1803,1674,1784,1402,1838,450,350,1102,705,1699,1631,1785,405,480,1315,1519,1305,1139,363,844,334,962,1126,1288,1014,506,831,1619,1121,554,1371,749,108,476,1361,984,368,376,234,321,1542,1165,1772,1177,702,1309,939,1908,1470,1989,1835,1717,1001,276,1763,180,298,25,988,1615,987,713,1250,463,1691,855,243,690,1055,1562,958,636,426,1012,1185,622,671,203,1742,1694,801,712,605,744,264,1665,1510,517,1464,42,1257,852,1185,1046,1739,1589,1193,1174,1772,1893,1408,960,1815,793,1897,1766,690,1928,1154,267,1434,145,555,970,1654,79,1907,1658,763,22,961,656,346,1879,79,300,530,341,421,325,1017,1159,279,1703,885,130,359,1501,1777,1800,1765,666,180,1179,1953,717,976,321,975,1957,655,1714,1942,55,1355,477,1524,1691,1540,1699,743,1865,1887,439,943,1017,816,1465,830,164,1605,677,869,2029,199,1224,1431,56,1868,294,384,1609,533,190,1932,469,1323,616,608,1253,201,1141,1466,398,1999,863,286,625,1096,724,167,2003,689,537,48,1489,1636,335,733,1146,1196,1559,1485,13,1040,281,1087,1187,1085,1010,165,1351,1239,978,1998,905,1927,1709,1756,219,551,1501,843,871,398,1557,1806,949,1962,557,1035,993,968,1771,463,2011,575,1128,1736,81,1779,1620,183,1232,301,565,339,361,1205,1167,1604,444,1831,1493,1986,1815,466,1971,914,1809,211,1159,1810,543,493,242,1605,945,1088,565,631,1168,259,1462,1852,908,1365,1259,1710,238,1367,108,1440,16,1817,1994,187,1425,858,1806,1420,455,256,1395,1369,959,1284,1503,287,1175,694,264,1362,86,1205,1826,870,1729,642,552,1190,321,1110,974,1974,1980,114,1360,1739,429,1705,208,1394,723,1183,1572,1971,1090,1786,1868,448,1825,933,47,1813,773,1529,1197,1707,1217,301,2031,982,1726,1474,1655,752,1309,1290,1212,917,1359,1969,1898,573,1175,875,1986,560,459,74,1612,991,1070,1445,490,321,1286,1170,1484,590,828,741,6,318,616,1658,707,1074,578,1594,1162,1029,850,950,1816,970,1019,1013,533,400,1829,1740,1876,1455,1266,822,998,1825,177,598,1851,460,1800,345,2044,1344,1735,362,910,1321,736,1585,2034,418,1434,1498,1143,1931,1513,1690,1028,1507,1914,1529,1523,157,367,805,1817,159,1606,1296,157,1961,727,1565,1152,507,305,1815,924,1125,1589,1755,1532,162,364,217,1522,1101,410,1106,718,1986,1264,1848,818,2,2027,1620,485,1908,661,1264,1458,726,809,910,1349,832,602,1675,1053,1428,435,599,2016,618,1352,81,251,1225,1114,1387,1410,1632,1141,256,1084,1814,1852,1282,10,1633,1316,896,612,638,1810,1594,1629,1425,1916,513,662,688,1187,504,1441,1819,187,699,935,1469,1498,1004,1561,805,824,94,1651,474,1630,1398,564,1294,1289,2040,1749,220,1785,243,878,1521,1315,364,30,442,1887,244,416,1560,1047,1944,1573,1437,782,1690,187,500,797,281,249,250,974,146,1150,1068,225,718,2010,288,1311,1845,412,1050,520,322,1160,984,1900,1982,1938,1312,171,1372,328,443,316,838,1876,1975,1143,1732,362,1905,744,1941,1508,1948,0),
   (0,0,0,0,-1,0,-1,0,0,0,1,0,0,0,0,0,0,-1,0,0,0,1,1,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,-1,0,0,0,-1,-1,0,0,0,0,0,0,0,0,1,0,0,0,0,0,1,1,0,-1,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,1,1,0,0,0,0,0,0,0,-1,0,0,0,0,1,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,-1,0,0,1,0,0,0,0,0,0,0,1,0,-1,0,0,0,0,0,0,0,0,0,-1,0,0,0,-1,0,0,0,1,0,0,0,0,0,0,0,0,1,0,0,0,0,-1,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,-1,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,0,0,0,1,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,1,0,0,0,1,0,0,0,0,0,-1,1,0,0,0,0,0,0,0,-1,-1,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,-1,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,-1,0,-1,0,0,0,0,0,0,1,0,1,0,0,-1,0,0,0,0,0,-1,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,1,0,0,-1,1,0,1,0,0,0,-1,0,0,1,0,-1,-1,0,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,0,-1,0,0,0,0,0,0,0,0,0,1,0,-1,0,1,0,0,0,0,0,0,-1,-1,1,0,0,0,0,0,0,0,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,0,0,0,0,0,1,-1,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,-1,0,0,1,0,0,0,0,0,0,0,0,0,0,-1,-1,0,0,0,-1,0,1,0,-1,0,0,0,0,0,0,0,0,0,0,0,0,-1,0,0,1,0,0,0,0,0,0,0,0,0,0,-1,0,0,0,-1,0,0,0,-1,0,0,0,0,0,0,0,0,0,-1,0,0,0,0,0,0,-1,0,0,0,-1,0,0,0,0,0,0,0,1,0,1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,1,0,0,0,1,0,1,0,0,0,0,-1,0,-1,0,1,0,0),
   '1',
   (486, 251, 2019, 423, 1295, 1109, 1045, 1240, 366, 353, 1411, 1238, 1126, 1145, 362, 1101, 2022, 1173, 270, 238, 588, 580, 698, 951, 842, 1174, 508, 545, 852, 1539, 1571, 1834, 590, 1536, 1172, 1849, 1059, 918, 1194, 667, 993, 1163, 916, 107, 722, 1319, 1750, 1950, 808, 716, 1849, 1077, 1229, 691, 979, 245, 215, 121, 1943, 1839, 711, 209, 1964, 1533, 1852, 1612, 1021, 1839, 853, 1309, 1540, 1177, 936, 80, 284, 359, 1899, 377, 6, 1214, 794, 899, 1034, 926, 926, 1941, 1163, 1264, 1544, 1163, 1123, 994, 675, 1890, 132, 763, 830, 892, 669, 1608, 502, 1717, 1309, 1385, 394, 696, 763, 1636, 827, 1000, 708, 1437, 1131, 1351, 621, 1801, 1063, 706, 672, 1703, 1848, 2033, 540, 554, 1006, 1725, 1514, 843, 299, 2010, 614, 1143, 1766, 1185, 820, 185, 168, 1023, 579, 1649, 356, 1586, 1804, 84, 969, 518, 113, 1920, 1324, 615, 1976, 299, 189, 1402, 436, 1085, 1088, 1534, 1247, 550, 2012, 857, 1161, 1356, 172, 784, 1650, 522, 377, 433, 1741, 106, 1094, 10, 1685, 1666, 289, 1070, 751, 1715, 390, 771, 590, 807, 1173, 596, 441, 239, 322, 1023, 991, 232, 770, 1529, 229, 283, 962, 70, 1830, 1261, 1515, 1756, 386, 1268, 1528, 458, 383, 1119, 133, 113, 703, 1848, 769, 536, 1588, 1355, 305, 928, 696, 766, 324, 237, 1786, 2025, 1227, 383, 1511, 1504, 1973, 1730, 1845, 991, 920, 966, 211, 844, 1726, 1394, 1618, 1100, 1086, 1782, 1365, 1304, 1029, 1593, 716, 1693, 694, 1143, 1365, 1667, 1801, 673, 1941, 1781, 1050, 525, 355, 1407, 1681, 66, 1997, 1898, 1160, 493, 1503, 808, 978, 356, 993, 81, 6, 1305, 704, 536, 1947, 1970, 445, 1614, 1745, 256, 417, 1190, 693, 1496, 847, 1490, 1529, 134, 997, 1127, 629, 1466, 409, 1786, 173, 1999, 289, 66, 168, 1003, 1688, 47, 1715, 1439, 716, 1231, 1817, 1777, 1905, 736, 681, 188, 1251, 448, 89, 706, 1961, 2014, 604, 1187, 1649, 836, 1223, 336, 172, 858, 2016, 2017, 351, 37, 2027, 1280, 109, 1115, 1043, 1335, 454, 17, 1665, 1501, 1363, 1151, 1522, 2022, 304, 882, 2011, 425, 1136, 73, 90, 1930, 999, 998, 1340, 669, 52, 714, 1922, 1646, 1561, 1142, 145, 1971, 1544, 1571, 842, 1413, 1670, 1641, 1847, 216, 814, 1, 1259, 637, 115, 1542, 2036, 1818, 9, 1311, 1233, 1903, 371, 1686, 1642, 72, 1336, 414, 1626, 1656, 539, 835, 144, 1629, 993, 1117, 1829, 1266, 1094, 379, 2012, 799, 2041, 59, 2027, 1450, 618, 110, 1756, 398, 408, 1783, 873, 1970, 1030, 1177, 1916, 1643, 1079, 1816, 609, 1560, 258, 1303, 1164, 1126, 828, 1108, 164, 908, 995, 1000, 179, 1087, 1682, 1479, 2018, 1015, 561, 1143, 3, 1506, 677, 565, 478, 837, 205, 324, 277, 864, 1368, 348, 1085, 1302, 1516, 136, 445, 547, 655, 271, 423, 778, 1136, 802, 1995, 1890, 1708, 1104, 1263, 1696, 482, 1025, 818, 1619, 1264, 1065, 1930, 1128, 524, 643, 1933, 953, 276, 1101, 1053, 1303, 1010, 1047, 209, 383, 491, 215, 492, 1164, 30, 813, 1392, 770, 341, 1945, 1935, 776, 869, 1973, 189, 2025, 1422, 1626, 1184, 1103, 4, 1905, 1288, 1832, 1977, 1004, 1604, 614, 532, 769, 1609, 1528, 829, 1505, 490, 1638, 1656, 1270, 1717, 374, 316, 862, 1302, 120, 1280, 1599, 1487, 101, 1708, 889, 735, 1662, 1412, 998, 506, 1082, 1391, 1468, 493, 974, 1600, 168, 972, 1989, 1169, 704, 650, 2030, 900, 1285, 51, 1753, 747, 1612, 180, 57, 953, 1215, 252, 127, 280, 780, 1653, 223, 1761, 1220, 568, 1574, 356, 6, 58, 1382, 566, 512, 212, 636, 1621, 270, 1894, 467, 1214, 1350, 1157, 1515, 1325, 1893, 1135, 568, 1970, 296, 1781, 900, 1952, 297, 541, 887, 1636, 424, 767, 1443, 945, 1560, 574, 1145, 0)
   );
end process;   
   
end a1;